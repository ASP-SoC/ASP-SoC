-------------------------------------------------------------------------------
-- Title      : Testbench Signal Delay Left and Right
-------------------------------------------------------------------------------
-- File       : tbDelay-Bhv-ea.vhd
-- Author     : Michael Wurm
-------------------------------------------------------------------------------
-- Description: Testbench, tests basic functions of unit Delay
-------------------------------------------------------------------------------
-- Copyright (c) 2017 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author    Description
-- 2017-06-06  1.0      MikeW     Created
-------------------------------------------------------------------------------


entity tbDelay is
end entity tbDelay;

architecture bhv of tbDelay is

begin


end architecture bhv;
