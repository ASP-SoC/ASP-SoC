-------------------------------------------------------------------------------
-- Title      : Equalizer Project Package
-------------------------------------------------------------------------------
-- Description: Type definitions and filter coefficients for unit Equalizer
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ieee_proposed;
use ieee_proposed.fixed_pkg.all;
use ieee_proposed.fixed_float_types.all;

package PkgEqualizer is

  constant cNumOfBands       : natural :=  10;
  constant cFilterCoeffWidth : natural :=  24;
  constant cEQBandpassOrder  : natural :=  79;

  subtype aFilterCoeff is u_sfixed(0 downto -(cFilterCoeffWidth-1));
  type aMemory is array (natural range <>) of aFilterCoeff;

  subtype fract_real is real range
    -1.0 to 0.99999999999999999999999999999999999999999999999999999999999999999;
  type aCoeffMemory is array (natural range <>) of fract_real;
  type aEQBandpassSet is array(natural range<>) of aCoeffMemory(0 to cEQBandpassOrder);

  constant cCoeffBandpass0 : aCoeffMemory(0 to cEQBandpassOrder) := (
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9
    );
  constant cCoeffBandpass1 : aCoeffMemory(0 to cEQBandpassOrder) := (
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9
  );
  constant cCoeffBandpass2 : aCoeffMemory(0 to cEQBandpassOrder) := (
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9
  );
  constant cCoeffBandpass3 : aCoeffMemory(0 to cEQBandpassOrder) := (
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9
  );
  constant cCoeffBandpass4 : aCoeffMemory(0 to cEQBandpassOrder) := (
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9
  );
  constant cCoeffBandpass5 : aCoeffMemory(0 to cEQBandpassOrder) := (
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9
  );
  constant cCoeffBandpass6 : aCoeffMemory(0 to cEQBandpassOrder) := (
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9
  );
  constant cCoeffBandpass7 : aCoeffMemory(0 to cEQBandpassOrder) := (
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9
  );
  constant cCoeffBandpass8 : aCoeffMemory(0 to cEQBandpassOrder) := (
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9
  );
  constant cCoeffBandpass9 : aCoeffMemory(0 to cEQBandpassOrder) := (
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,
    0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9,0.9
  );

  ------------------------------------------------------------------------------
  -- Function Definitions
  ------------------------------------------------------------------------------
  function ResizeTruncAbsVal (
    arg      : u_sfixed;  -- input
    size_res : u_sfixed)  -- for size only
    return sfixed;

end PkgEqualizer;

package body PkgEqualizer is

  function ResizeTruncAbsVal (
    arg : u_sfixed;
    size_res : u_sfixed)
  return sfixed is
    variable lsb : u_sfixed(size_res'range) := (others => '0');
    variable tmp : u_sfixed(size_res'high+1 downto size_res'low) := (others => '0');
  begin
    lsb(lsb'low) := '1';
    tmp(size_res'range) := resize(arg => arg,
                           left_index => size_res'high,
                           right_index => size_res'low,
                           round_style => fixed_truncate,
                           overflow_style => fixed_saturate);

    if tmp < 0 and arg > -1 then
      tmp := tmp(size_res'range) + lsb;
    end if;
    return tmp(size_res'range);
  end function ResizeTruncAbsVal;

end PkgEqualizer;
