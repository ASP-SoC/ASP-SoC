architecture Struct of PlatformHps is

begin  -- architecture Struct

  

end architecture Struct;
