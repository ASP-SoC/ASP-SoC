architecture Struct of AudioSignalProcessingBlock is

begin  -- architecture Struct



end architecture Struct;
