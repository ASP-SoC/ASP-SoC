library ieee;
use ieee.std_logic_1164.all;

use work.Global.all;

package sin_4096 is

  -- sin table with 4096 values
  constant sin_table_c : fract_set_t := (
    0.00076699, 0.00230097, 0.00383494, 0.00536891, 0.00690286, 0.00843679, 0.00997071, 0.01150460, 0.01303847, 0.01457230,
    0.01610610, 0.01763986, 0.01917358, 0.02070726, 0.02224089, 0.02377446, 0.02530798, 0.02684144, 0.02837484, 0.02990816,
    0.03144142, 0.03297461, 0.03450772, 0.03604074, 0.03757368, 0.03910654, 0.04063930, 0.04217196, 0.04370453, 0.04523699,
    0.04676935, 0.04830159, 0.04983373, 0.05136574, 0.05289764, 0.05442941, 0.05596105, 0.05749256, 0.05902393, 0.06055517,
    0.06208627, 0.06361721, 0.06514801, 0.06667866, 0.06820914, 0.06973947, 0.07126963, 0.07279963, 0.07432945, 0.07585910,
    0.07738857, 0.07891786, 0.08044697, 0.08197588, 0.08350460, 0.08503312, 0.08656145, 0.08808957, 0.08961748, 0.09114519,
    0.09267267, 0.09419994, 0.09572699, 0.09725381, 0.09878041, 0.10030677, 0.10183290, 0.10335878, 0.10488442, 0.10640982,
    0.10793497, 0.10945986, 0.11098449, 0.11250886, 0.11403297, 0.11555681, 0.11708038, 0.11860367, 0.12012669, 0.12164942,
    0.12317186, 0.12469402, 0.12621588, 0.12773744, 0.12925870, 0.13077966, 0.13230032, 0.13382066, 0.13534068, 0.13686039,
    0.13837977, 0.13989883, 0.14141756, 0.14293596, 0.14445402, 0.14597174, 0.14748912, 0.14900615, 0.15052283, 0.15203916,
    0.15355512, 0.15507073, 0.15658597, 0.15810085, 0.15961535, 0.16112947, 0.16264322, 0.16415658, 0.16566956, 0.16718215,
    0.16869434, 0.17020614, 0.17171754, 0.17322853, 0.17473911, 0.17624929, 0.17775905, 0.17926839, 0.18077731, 0.18228580,
    0.18379387, 0.18530150, 0.18680870, 0.18831545, 0.18982177, 0.19132763, 0.19283305, 0.19433801, 0.19584252, 0.19734656,
    0.19885014, 0.20035326, 0.20185590, 0.20335806, 0.20485975, 0.20636096, 0.20786168, 0.20936191, 0.21086164, 0.21236089,
    0.21385963, 0.21535787, 0.21685560, 0.21835282, 0.21984953, 0.22134572, 0.22284139, 0.22433654, 0.22583115, 0.22732524,
    0.22881879, 0.23031180, 0.23180428, 0.23329620, 0.23478758, 0.23627840, 0.23776867, 0.23925838, 0.24074752, 0.24223610,
    0.24372411, 0.24521155, 0.24669841, 0.24818469, 0.24967038, 0.25115549, 0.25264000, 0.25412392, 0.25560725, 0.25708997,
    0.25857208, 0.26005359, 0.26153449, 0.26301477, 0.26449443, 0.26597347, 0.26745189, 0.26892967, 0.27040682, 0.27188334,
    0.27335921, 0.27483445, 0.27630903, 0.27778297, 0.27925625, 0.28072887, 0.28220084, 0.28367214, 0.28514277, 0.28661273,
    0.28808202, 0.28955063, 0.29101856, 0.29248580, 0.29395235, 0.29541822, 0.29688339, 0.29834785, 0.29981162, 0.30127468,
    0.30273704, 0.30419868, 0.30565960, 0.30711981, 0.30857929, 0.31003805, 0.31149607, 0.31295337, 0.31440993, 0.31586575,
    0.31732082, 0.31877515, 0.32022873, 0.32168155, 0.32313362, 0.32458492, 0.32603547, 0.32748524, 0.32893425, 0.33038248,
    0.33182994, 0.33327661, 0.33472250, 0.33616760, 0.33761191, 0.33905543, 0.34049814, 0.34194006, 0.34338117, 0.34482148,
    0.34626097, 0.34769965, 0.34913751, 0.35057455, 0.35201076, 0.35344614, 0.35488070, 0.35631442, 0.35774730, 0.35917933,
    0.36061053, 0.36204087, 0.36347036, 0.36489900, 0.36632678, 0.36775370, 0.36917975, 0.37060493, 0.37202924, 0.37345267,
    0.37487523, 0.37629691, 0.37771769, 0.37913759, 0.38055660, 0.38197471, 0.38339193, 0.38480824, 0.38622364, 0.38763814,
    0.38905172, 0.39046439, 0.39187614, 0.39328697, 0.39469688, 0.39610585, 0.39751389, 0.39892100, 0.40032717, 0.40173239,
    0.40313667, 0.40454000, 0.40594238, 0.40734381, 0.40874428, 0.41014378, 0.41154232, 0.41293989, 0.41433649, 0.41573211,
    0.41712676, 0.41852043, 0.41991310, 0.42130480, 0.42269550, 0.42408520, 0.42547391, 0.42686162, 0.42824832, 0.42963401,
    0.43101870, 0.43240237, 0.43378502, 0.43516665, 0.43654726, 0.43792683, 0.43930538, 0.44068290, 0.44205938, 0.44343482,
    0.44480921, 0.44618256, 0.44755486, 0.44892610, 0.45029629, 0.45166542, 0.45303349, 0.45440049, 0.45576642, 0.45713128,
    0.45849506, 0.45985776, 0.46121939, 0.46257992, 0.46393937, 0.46529773, 0.46665499, 0.46801115, 0.46936622, 0.47072017,
    0.47207302, 0.47342476, 0.47477539, 0.47612490, 0.47747328, 0.47882055, 0.48016669, 0.48151169, 0.48285557, 0.48419831,
    0.48553990, 0.48688036, 0.48821967, 0.48955783, 0.49089484, 0.49223070, 0.49356540, 0.49489893, 0.49623130, 0.49756250,
    0.49889254, 0.50022139, 0.50154908, 0.50287558, 0.50420089, 0.50552503, 0.50684797, 0.50816972, 0.50949027, 0.51080962,
    0.51212778, 0.51344472, 0.51476046, 0.51607499, 0.51738830, 0.51870040, 0.52001128, 0.52132093, 0.52262935, 0.52393655,
    0.52524251, 0.52654724, 0.52785072, 0.52915297, 0.53045397, 0.53175372, 0.53305222, 0.53434947, 0.53564546, 0.53694019,
    0.53823365, 0.53952585, 0.54081678, 0.54210643, 0.54339482, 0.54468192, 0.54596774, 0.54725227, 0.54853552, 0.54981748,
    0.55109814, 0.55237751, 0.55365558, 0.55493234, 0.55620780, 0.55748195, 0.55875479, 0.56002631, 0.56129651, 0.56256540,
    0.56383296, 0.56509919, 0.56636410, 0.56762767, 0.56888990, 0.57015080, 0.57141036, 0.57266857, 0.57392543, 0.57518094,
    0.57643510, 0.57768790, 0.57893935, 0.58018943, 0.58143815, 0.58268549, 0.58393147, 0.58517607, 0.58641930, 0.58766114,
    0.58890161, 0.59014068, 0.59137837, 0.59261467, 0.59384957, 0.59508308, 0.59631518, 0.59754588, 0.59877518, 0.60000307,
    0.60122954, 0.60245460, 0.60367824, 0.60490046, 0.60612126, 0.60734063, 0.60855858, 0.60977509, 0.61099016, 0.61220380,
    0.61341600, 0.61462676, 0.61583606, 0.61704392, 0.61825033, 0.61945528, 0.62065878, 0.62186081, 0.62306138, 0.62426049,
    0.62545812, 0.62665429, 0.62784898, 0.62904219, 0.63023392, 0.63142417, 0.63261293, 0.63380021, 0.63498599, 0.63617028,
    0.63735307, 0.63853436, 0.63971415, 0.64089244, 0.64206921, 0.64324448, 0.64441823, 0.64559046, 0.64676118, 0.64793038,
    0.64909805, 0.65026419, 0.65142880, 0.65259188, 0.65375342, 0.65491343, 0.65607189, 0.65722881, 0.65838419, 0.65953801,
    0.66069028, 0.66184100, 0.66299016, 0.66413776, 0.66528380, 0.66642827, 0.66757118, 0.66871251, 0.66985227, 0.67099045,
    0.67212706, 0.67326208, 0.67439552, 0.67552737, 0.67665764, 0.67778631, 0.67891338, 0.68003886, 0.68116274, 0.68228501,
    0.68340568, 0.68452474, 0.68564219, 0.68675803, 0.68787225, 0.68898485, 0.69009583, 0.69120519, 0.69231292, 0.69341902,
    0.69452349, 0.69562633, 0.69672753, 0.69782709, 0.69892500, 0.70002128, 0.70111590, 0.70220888, 0.70330020, 0.70438987,
    0.70547788, 0.70656423, 0.70764892, 0.70873194, 0.70981330, 0.71089298, 0.71197099, 0.71304733, 0.71412199, 0.71519497,
    0.71626626, 0.71733587, 0.71840380, 0.71947003, 0.72053457, 0.72159741, 0.72265855, 0.72371800, 0.72477574, 0.72583178,
    0.72688611, 0.72793872, 0.72898963, 0.73003882, 0.73108629, 0.73213204, 0.73317607, 0.73421837, 0.73525895, 0.73629780,
    0.73733491, 0.73837029, 0.73940393, 0.74043583, 0.74146599, 0.74249440, 0.74352107, 0.74454598, 0.74556915, 0.74659056,
    0.74761021, 0.74862811, 0.74964424, 0.75065861, 0.75167121, 0.75268205, 0.75369111, 0.75469840, 0.75570391, 0.75670765,
    0.75770960, 0.75870977, 0.75970816, 0.76070476, 0.76169957, 0.76269258, 0.76368380, 0.76467323, 0.76566085, 0.76664668,
    0.76763070, 0.76861291, 0.76959331, 0.77057191, 0.77154869, 0.77252365, 0.77349680, 0.77446813, 0.77543763, 0.77640531,
    0.77737116, 0.77833519, 0.77929738, 0.78025774, 0.78121626, 0.78217294, 0.78312779, 0.78408079, 0.78503194, 0.78598125,
    0.78692871, 0.78787432, 0.78881807, 0.78975997, 0.79070001, 0.79163819, 0.79257450, 0.79350895, 0.79444154, 0.79537225,
    0.79630109, 0.79722806, 0.79815315, 0.79907637, 0.79999770, 0.80091715, 0.80183472, 0.80275040, 0.80366419, 0.80457609,
    0.80548610, 0.80639421, 0.80730042, 0.80820474, 0.80910715, 0.81000766, 0.81090626, 0.81180296, 0.81269774, 0.81359061,
    0.81448157, 0.81537061, 0.81625773, 0.81714293, 0.81802621, 0.81890757, 0.81978699, 0.82066449, 0.82154006, 0.82241369,
    0.82328539, 0.82415515, 0.82502297, 0.82588885, 0.82675279, 0.82761478, 0.82847482, 0.82933292, 0.83018906, 0.83104325,
    0.83189548, 0.83274576, 0.83359408, 0.83444043, 0.83528483, 0.83612725, 0.83696771, 0.83780620, 0.83864272, 0.83947726,
    0.84030983, 0.84114042, 0.84196904, 0.84279567, 0.84362032, 0.84444298, 0.84526365, 0.84608234, 0.84689904, 0.84771374,
    0.84852645, 0.84933716, 0.85014587, 0.85095259, 0.85175730, 0.85256000, 0.85336070, 0.85415940, 0.85495608, 0.85575075,
    0.85654340, 0.85733405, 0.85812267, 0.85890927, 0.85969386, 0.86047642, 0.86125695, 0.86203546, 0.86281194, 0.86358639,
    0.86435881, 0.86512920, 0.86589754, 0.86666385, 0.86742813, 0.86819036, 0.86895054, 0.86970869, 0.87046478, 0.87121883,
    0.87197083, 0.87272078, 0.87346867, 0.87421451, 0.87495829, 0.87570001, 0.87643967, 0.87717727, 0.87791280, 0.87864627,
    0.87937767, 0.88010700, 0.88083426, 0.88155945, 0.88228256, 0.88300360, 0.88372256, 0.88443944, 0.88515424, 0.88586695,
    0.88657759, 0.88728613, 0.88799259, 0.88869696, 0.88939923, 0.89009942, 0.89079751, 0.89149350, 0.89218739, 0.89287919,
    0.89356889, 0.89425648, 0.89494197, 0.89562535, 0.89630662, 0.89698579, 0.89766284, 0.89833779, 0.89901062, 0.89968133,
    0.90034993, 0.90101640, 0.90168076, 0.90234300, 0.90300311, 0.90366110, 0.90431696, 0.90497069, 0.90562229, 0.90627177,
    0.90691911, 0.90756431, 0.90820738, 0.90884832, 0.90948711, 0.91012377, 0.91075828, 0.91139065, 0.91202088, 0.91264896,
    0.91327489, 0.91389867, 0.91452030, 0.91513978, 0.91575711, 0.91637228, 0.91698530, 0.91759616, 0.91820486, 0.91881139,
    0.91941577, 0.92001798, 0.92061803, 0.92121591, 0.92181163, 0.92240517, 0.92299654, 0.92358575, 0.92417278, 0.92475763,
    0.92534031, 0.92592081, 0.92649913, 0.92707527, 0.92764923, 0.92822101, 0.92879060, 0.92935801, 0.92992323, 0.93048627,
    0.93104711, 0.93160576, 0.93216222, 0.93271649, 0.93326856, 0.93381844, 0.93436611, 0.93491159, 0.93545487, 0.93599595,
    0.93653483, 0.93707150, 0.93760597, 0.93813823, 0.93866828, 0.93919613, 0.93972176, 0.94024519, 0.94076640, 0.94128540,
    0.94180218, 0.94231675, 0.94282909, 0.94333923, 0.94384714, 0.94435283, 0.94485629, 0.94535754, 0.94585656, 0.94635335,
    0.94684792, 0.94734026, 0.94783037, 0.94831825, 0.94880389, 0.94928731, 0.94976849, 0.95024744, 0.95072415, 0.95119862,
    0.95167086, 0.95214085, 0.95260861, 0.95307412, 0.95353740, 0.95399842, 0.95445721, 0.95491374, 0.95536803, 0.95582007,
    0.95626987, 0.95671741, 0.95716270, 0.95760574, 0.95804652, 0.95848506, 0.95892133, 0.95935535, 0.95978711, 0.96021662,
    0.96064386, 0.96106884, 0.96149156, 0.96191202, 0.96233022, 0.96274615, 0.96315982, 0.96357122, 0.96398035, 0.96438721,
    0.96479181, 0.96519413, 0.96559418, 0.96599197, 0.96638747, 0.96678071, 0.96717167, 0.96756035, 0.96794676, 0.96833088,
    0.96871273, 0.96909231, 0.96946960, 0.96984460, 0.97021733, 0.97058778, 0.97095594, 0.97132181, 0.97168540, 0.97204670,
    0.97240572, 0.97276245, 0.97311689, 0.97346903, 0.97381889, 0.97416646, 0.97451173, 0.97485471, 0.97519540, 0.97553379,
    0.97586989, 0.97620369, 0.97653520, 0.97686440, 0.97719131, 0.97751592, 0.97783822, 0.97815823, 0.97847594, 0.97879134,
    0.97910444, 0.97941523, 0.97972372, 0.98002991, 0.98033379, 0.98063536, 0.98093462, 0.98123158, 0.98152623, 0.98181857,
    0.98210859, 0.98239631, 0.98268172, 0.98296481, 0.98324559, 0.98352405, 0.98380021, 0.98407404, 0.98434556, 0.98461477,
    0.98488166, 0.98514623, 0.98540848, 0.98566841, 0.98592603, 0.98618132, 0.98643429, 0.98668495, 0.98693328, 0.98717929,
    0.98742297, 0.98766433, 0.98790337, 0.98814008, 0.98837447, 0.98860653, 0.98883627, 0.98906368, 0.98928876, 0.98951151,
    0.98973194, 0.98995004, 0.99016580, 0.99037924, 0.99059035, 0.99079912, 0.99100557, 0.99120968, 0.99141146, 0.99161091,
    0.99180802, 0.99200280, 0.99219524, 0.99238535, 0.99257313, 0.99275857, 0.99294167, 0.99312244, 0.99330087, 0.99347697,
    0.99365072, 0.99382214, 0.99399122, 0.99415796, 0.99432236, 0.99448442, 0.99464414, 0.99480152, 0.99495656, 0.99510926,
    0.99525961, 0.99540763, 0.99555330, 0.99569663, 0.99583761, 0.99597626, 0.99611256, 0.99624651, 0.99637812, 0.99650739,
    0.99663431, 0.99675889, 0.99688112, 0.99700101, 0.99711855, 0.99723374, 0.99734659, 0.99745709, 0.99756524, 0.99767104,
    0.99777450, 0.99787561, 0.99797437, 0.99807079, 0.99816485, 0.99825657, 0.99834593, 0.99843295, 0.99851762, 0.99859994,
    0.99867991, 0.99875753, 0.99883280, 0.99890572, 0.99897628, 0.99904450, 0.99911037, 0.99917388, 0.99923505, 0.99929386,
    0.99935032, 0.99940443, 0.99945619, 0.99950560, 0.99955265, 0.99959735, 0.99963970, 0.99967970, 0.99971735, 0.99975264,
    0.99978558, 0.99981617, 0.99984441, 0.99987029, 0.99989382, 0.99991500, 0.99993382, 0.99995029, 0.99996441, 0.99997617,
    0.99998559, 0.99999265, 0.99999735, 0.99999971, 0.99999971, 0.99999735, 0.99999265, 0.99998559, 0.99997617, 0.99996441,
    0.99995029, 0.99993382, 0.99991500, 0.99989382, 0.99987029, 0.99984441, 0.99981617, 0.99978558, 0.99975264, 0.99971735,
    0.99967970, 0.99963970, 0.99959735, 0.99955265, 0.99950560, 0.99945619, 0.99940443, 0.99935032, 0.99929386, 0.99923505,
    0.99917388, 0.99911037, 0.99904450, 0.99897628, 0.99890572, 0.99883280, 0.99875753, 0.99867991, 0.99859994, 0.99851762,
    0.99843295, 0.99834593, 0.99825657, 0.99816485, 0.99807079, 0.99797437, 0.99787561, 0.99777450, 0.99767104, 0.99756524,
    0.99745709, 0.99734659, 0.99723374, 0.99711855, 0.99700101, 0.99688112, 0.99675889, 0.99663431, 0.99650739, 0.99637812,
    0.99624651, 0.99611256, 0.99597626, 0.99583761, 0.99569663, 0.99555330, 0.99540763, 0.99525961, 0.99510926, 0.99495656,
    0.99480152, 0.99464414, 0.99448442, 0.99432236, 0.99415796, 0.99399122, 0.99382214, 0.99365072, 0.99347697, 0.99330087,
    0.99312244, 0.99294167, 0.99275857, 0.99257313, 0.99238535, 0.99219524, 0.99200280, 0.99180802, 0.99161091, 0.99141146,
    0.99120968, 0.99100557, 0.99079912, 0.99059035, 0.99037924, 0.99016580, 0.98995004, 0.98973194, 0.98951151, 0.98928876,
    0.98906368, 0.98883627, 0.98860653, 0.98837447, 0.98814008, 0.98790337, 0.98766433, 0.98742297, 0.98717929, 0.98693328,
    0.98668495, 0.98643429, 0.98618132, 0.98592603, 0.98566841, 0.98540848, 0.98514623, 0.98488166, 0.98461477, 0.98434556,
    0.98407404, 0.98380021, 0.98352405, 0.98324559, 0.98296481, 0.98268172, 0.98239631, 0.98210859, 0.98181857, 0.98152623,
    0.98123158, 0.98093462, 0.98063536, 0.98033379, 0.98002991, 0.97972372, 0.97941523, 0.97910444, 0.97879134, 0.97847594,
    0.97815823, 0.97783822, 0.97751592, 0.97719131, 0.97686440, 0.97653520, 0.97620369, 0.97586989, 0.97553379, 0.97519540,
    0.97485471, 0.97451173, 0.97416646, 0.97381889, 0.97346903, 0.97311689, 0.97276245, 0.97240572, 0.97204670, 0.97168540,
    0.97132181, 0.97095594, 0.97058778, 0.97021733, 0.96984460, 0.96946960, 0.96909231, 0.96871273, 0.96833088, 0.96794676,
    0.96756035, 0.96717167, 0.96678071, 0.96638747, 0.96599197, 0.96559418, 0.96519413, 0.96479181, 0.96438721, 0.96398035,
    0.96357122, 0.96315982, 0.96274615, 0.96233022, 0.96191202, 0.96149156, 0.96106884, 0.96064386, 0.96021662, 0.95978711,
    0.95935535, 0.95892133, 0.95848506, 0.95804652, 0.95760574, 0.95716270, 0.95671741, 0.95626987, 0.95582007, 0.95536803,
    0.95491374, 0.95445721, 0.95399842, 0.95353740, 0.95307412, 0.95260861, 0.95214085, 0.95167086, 0.95119862, 0.95072415,
    0.95024744, 0.94976849, 0.94928731, 0.94880389, 0.94831825, 0.94783037, 0.94734026, 0.94684792, 0.94635335, 0.94585656,
    0.94535754, 0.94485629, 0.94435283, 0.94384714, 0.94333923, 0.94282909, 0.94231675, 0.94180218, 0.94128540, 0.94076640,
    0.94024519, 0.93972176, 0.93919613, 0.93866828, 0.93813823, 0.93760597, 0.93707150, 0.93653483, 0.93599595, 0.93545487,
    0.93491159, 0.93436611, 0.93381844, 0.93326856, 0.93271649, 0.93216222, 0.93160576, 0.93104711, 0.93048627, 0.92992323,
    0.92935801, 0.92879060, 0.92822101, 0.92764923, 0.92707527, 0.92649913, 0.92592081, 0.92534031, 0.92475763, 0.92417278,
    0.92358575, 0.92299654, 0.92240517, 0.92181163, 0.92121591, 0.92061803, 0.92001798, 0.91941577, 0.91881139, 0.91820486,
    0.91759616, 0.91698530, 0.91637228, 0.91575711, 0.91513978, 0.91452030, 0.91389867, 0.91327489, 0.91264896, 0.91202088,
    0.91139065, 0.91075828, 0.91012377, 0.90948711, 0.90884832, 0.90820738, 0.90756431, 0.90691911, 0.90627177, 0.90562229,
    0.90497069, 0.90431696, 0.90366110, 0.90300311, 0.90234300, 0.90168076, 0.90101640, 0.90034993, 0.89968133, 0.89901062,
    0.89833779, 0.89766284, 0.89698579, 0.89630662, 0.89562535, 0.89494197, 0.89425648, 0.89356889, 0.89287919, 0.89218739,
    0.89149350, 0.89079751, 0.89009942, 0.88939923, 0.88869696, 0.88799259, 0.88728613, 0.88657759, 0.88586695, 0.88515424,
    0.88443944, 0.88372256, 0.88300360, 0.88228256, 0.88155945, 0.88083426, 0.88010700, 0.87937767, 0.87864627, 0.87791280,
    0.87717727, 0.87643967, 0.87570001, 0.87495829, 0.87421451, 0.87346867, 0.87272078, 0.87197083, 0.87121883, 0.87046478,
    0.86970869, 0.86895054, 0.86819036, 0.86742813, 0.86666385, 0.86589754, 0.86512920, 0.86435881, 0.86358639, 0.86281194,
    0.86203546, 0.86125695, 0.86047642, 0.85969386, 0.85890927, 0.85812267, 0.85733405, 0.85654340, 0.85575075, 0.85495608,
    0.85415940, 0.85336070, 0.85256000, 0.85175730, 0.85095259, 0.85014587, 0.84933716, 0.84852645, 0.84771374, 0.84689904,
    0.84608234, 0.84526365, 0.84444298, 0.84362032, 0.84279567, 0.84196904, 0.84114042, 0.84030983, 0.83947726, 0.83864272,
    0.83780620, 0.83696771, 0.83612725, 0.83528483, 0.83444043, 0.83359408, 0.83274576, 0.83189548, 0.83104325, 0.83018906,
    0.82933292, 0.82847482, 0.82761478, 0.82675279, 0.82588885, 0.82502297, 0.82415515, 0.82328539, 0.82241369, 0.82154006,
    0.82066449, 0.81978699, 0.81890757, 0.81802621, 0.81714293, 0.81625773, 0.81537061, 0.81448157, 0.81359061, 0.81269774,
    0.81180296, 0.81090626, 0.81000766, 0.80910715, 0.80820474, 0.80730042, 0.80639421, 0.80548610, 0.80457609, 0.80366419,
    0.80275040, 0.80183472, 0.80091715, 0.79999770, 0.79907637, 0.79815315, 0.79722806, 0.79630109, 0.79537225, 0.79444154,
    0.79350895, 0.79257450, 0.79163819, 0.79070001, 0.78975997, 0.78881807, 0.78787432, 0.78692871, 0.78598125, 0.78503194,
    0.78408079, 0.78312779, 0.78217294, 0.78121626, 0.78025774, 0.77929738, 0.77833519, 0.77737116, 0.77640531, 0.77543763,
    0.77446813, 0.77349680, 0.77252365, 0.77154869, 0.77057191, 0.76959331, 0.76861291, 0.76763070, 0.76664668, 0.76566085,
    0.76467323, 0.76368380, 0.76269258, 0.76169957, 0.76070476, 0.75970816, 0.75870977, 0.75770960, 0.75670765, 0.75570391,
    0.75469840, 0.75369111, 0.75268205, 0.75167121, 0.75065861, 0.74964424, 0.74862811, 0.74761021, 0.74659056, 0.74556915,
    0.74454598, 0.74352107, 0.74249440, 0.74146599, 0.74043583, 0.73940393, 0.73837029, 0.73733491, 0.73629780, 0.73525895,
    0.73421837, 0.73317607, 0.73213204, 0.73108629, 0.73003882, 0.72898963, 0.72793872, 0.72688611, 0.72583178, 0.72477574,
    0.72371800, 0.72265855, 0.72159741, 0.72053457, 0.71947003, 0.71840380, 0.71733587, 0.71626626, 0.71519497, 0.71412199,
    0.71304733, 0.71197099, 0.71089298, 0.70981330, 0.70873194, 0.70764892, 0.70656423, 0.70547788, 0.70438987, 0.70330020,
    0.70220888, 0.70111590, 0.70002128, 0.69892500, 0.69782709, 0.69672753, 0.69562633, 0.69452349, 0.69341902, 0.69231292,
    0.69120519, 0.69009583, 0.68898485, 0.68787225, 0.68675803, 0.68564219, 0.68452474, 0.68340568, 0.68228501, 0.68116274,
    0.68003886, 0.67891338, 0.67778631, 0.67665764, 0.67552737, 0.67439552, 0.67326208, 0.67212706, 0.67099045, 0.66985227,
    0.66871251, 0.66757118, 0.66642827, 0.66528380, 0.66413776, 0.66299016, 0.66184100, 0.66069028, 0.65953801, 0.65838419,
    0.65722881, 0.65607189, 0.65491343, 0.65375342, 0.65259188, 0.65142880, 0.65026419, 0.64909805, 0.64793038, 0.64676118,
    0.64559046, 0.64441823, 0.64324448, 0.64206921, 0.64089244, 0.63971415, 0.63853436, 0.63735307, 0.63617028, 0.63498599,
    0.63380021, 0.63261293, 0.63142417, 0.63023392, 0.62904219, 0.62784898, 0.62665429, 0.62545812, 0.62426049, 0.62306138,
    0.62186081, 0.62065878, 0.61945528, 0.61825033, 0.61704392, 0.61583606, 0.61462676, 0.61341600, 0.61220380, 0.61099016,
    0.60977509, 0.60855858, 0.60734063, 0.60612126, 0.60490046, 0.60367824, 0.60245460, 0.60122954, 0.60000307, 0.59877518,
    0.59754588, 0.59631518, 0.59508308, 0.59384957, 0.59261467, 0.59137837, 0.59014068, 0.58890161, 0.58766114, 0.58641930,
    0.58517607, 0.58393147, 0.58268549, 0.58143815, 0.58018943, 0.57893935, 0.57768790, 0.57643510, 0.57518094, 0.57392543,
    0.57266857, 0.57141036, 0.57015080, 0.56888990, 0.56762767, 0.56636410, 0.56509919, 0.56383296, 0.56256540, 0.56129651,
    0.56002631, 0.55875479, 0.55748195, 0.55620780, 0.55493234, 0.55365558, 0.55237751, 0.55109814, 0.54981748, 0.54853552,
    0.54725227, 0.54596774, 0.54468192, 0.54339482, 0.54210643, 0.54081678, 0.53952585, 0.53823365, 0.53694019, 0.53564546,
    0.53434947, 0.53305222, 0.53175372, 0.53045397, 0.52915297, 0.52785072, 0.52654724, 0.52524251, 0.52393655, 0.52262935,
    0.52132093, 0.52001128, 0.51870040, 0.51738830, 0.51607499, 0.51476046, 0.51344472, 0.51212778, 0.51080962, 0.50949027,
    0.50816972, 0.50684797, 0.50552503, 0.50420089, 0.50287558, 0.50154908, 0.50022139, 0.49889254, 0.49756250, 0.49623130,
    0.49489893, 0.49356540, 0.49223070, 0.49089484, 0.48955783, 0.48821967, 0.48688036, 0.48553990, 0.48419831, 0.48285557,
    0.48151169, 0.48016669, 0.47882055, 0.47747328, 0.47612490, 0.47477539, 0.47342476, 0.47207302, 0.47072017, 0.46936622,
    0.46801115, 0.46665499, 0.46529773, 0.46393937, 0.46257992, 0.46121939, 0.45985776, 0.45849506, 0.45713128, 0.45576642,
    0.45440049, 0.45303349, 0.45166542, 0.45029629, 0.44892610, 0.44755486, 0.44618256, 0.44480921, 0.44343482, 0.44205938,
    0.44068290, 0.43930538, 0.43792683, 0.43654726, 0.43516665, 0.43378502, 0.43240237, 0.43101870, 0.42963401, 0.42824832,
    0.42686162, 0.42547391, 0.42408520, 0.42269550, 0.42130480, 0.41991310, 0.41852043, 0.41712676, 0.41573211, 0.41433649,
    0.41293989, 0.41154232, 0.41014378, 0.40874428, 0.40734381, 0.40594238, 0.40454000, 0.40313667, 0.40173239, 0.40032717,
    0.39892100, 0.39751389, 0.39610585, 0.39469688, 0.39328697, 0.39187614, 0.39046439, 0.38905172, 0.38763814, 0.38622364,
    0.38480824, 0.38339193, 0.38197471, 0.38055660, 0.37913759, 0.37771769, 0.37629691, 0.37487523, 0.37345267, 0.37202924,
    0.37060493, 0.36917975, 0.36775370, 0.36632678, 0.36489900, 0.36347036, 0.36204087, 0.36061053, 0.35917933, 0.35774730,
    0.35631442, 0.35488070, 0.35344614, 0.35201076, 0.35057455, 0.34913751, 0.34769965, 0.34626097, 0.34482148, 0.34338117,
    0.34194006, 0.34049814, 0.33905543, 0.33761191, 0.33616760, 0.33472250, 0.33327661, 0.33182994, 0.33038248, 0.32893425,
    0.32748524, 0.32603547, 0.32458492, 0.32313362, 0.32168155, 0.32022873, 0.31877515, 0.31732082, 0.31586575, 0.31440993,
    0.31295337, 0.31149607, 0.31003805, 0.30857929, 0.30711981, 0.30565960, 0.30419868, 0.30273704, 0.30127468, 0.29981162,
    0.29834785, 0.29688339, 0.29541822, 0.29395235, 0.29248580, 0.29101856, 0.28955063, 0.28808202, 0.28661273, 0.28514277,
    0.28367214, 0.28220084, 0.28072887, 0.27925625, 0.27778297, 0.27630903, 0.27483445, 0.27335921, 0.27188334, 0.27040682,
    0.26892967, 0.26745189, 0.26597347, 0.26449443, 0.26301477, 0.26153449, 0.26005359, 0.25857208, 0.25708997, 0.25560725,
    0.25412392, 0.25264000, 0.25115549, 0.24967038, 0.24818469, 0.24669841, 0.24521155, 0.24372411, 0.24223610, 0.24074752,
    0.23925838, 0.23776867, 0.23627840, 0.23478758, 0.23329620, 0.23180428, 0.23031180, 0.22881879, 0.22732524, 0.22583115,
    0.22433654, 0.22284139, 0.22134572, 0.21984953, 0.21835282, 0.21685560, 0.21535787, 0.21385963, 0.21236089, 0.21086164,
    0.20936191, 0.20786168, 0.20636096, 0.20485975, 0.20335806, 0.20185590, 0.20035326, 0.19885014, 0.19734656, 0.19584252,
    0.19433801, 0.19283305, 0.19132763, 0.18982177, 0.18831545, 0.18680870, 0.18530150, 0.18379387, 0.18228580, 0.18077731,
    0.17926839, 0.17775905, 0.17624929, 0.17473911, 0.17322853, 0.17171754, 0.17020614, 0.16869434, 0.16718215, 0.16566956,
    0.16415658, 0.16264322, 0.16112947, 0.15961535, 0.15810085, 0.15658597, 0.15507073, 0.15355512, 0.15203916, 0.15052283,
    0.14900615, 0.14748912, 0.14597174, 0.14445402, 0.14293596, 0.14141756, 0.13989883, 0.13837977, 0.13686039, 0.13534068,
    0.13382066, 0.13230032, 0.13077966, 0.12925870, 0.12773744, 0.12621588, 0.12469402, 0.12317186, 0.12164942, 0.12012669,
    0.11860367, 0.11708038, 0.11555681, 0.11403297, 0.11250886, 0.11098449, 0.10945986, 0.10793497, 0.10640982, 0.10488442,
    0.10335878, 0.10183290, 0.10030677, 0.09878041, 0.09725381, 0.09572699, 0.09419994, 0.09267267, 0.09114519, 0.08961748,
    0.08808957, 0.08656145, 0.08503312, 0.08350460, 0.08197588, 0.08044697, 0.07891786, 0.07738857, 0.07585910, 0.07432945,
    0.07279963, 0.07126963, 0.06973947, 0.06820914, 0.06667866, 0.06514801, 0.06361721, 0.06208627, 0.06055517, 0.05902393,
    0.05749256, 0.05596105, 0.05442941, 0.05289764, 0.05136574, 0.04983373, 0.04830159, 0.04676935, 0.04523699, 0.04370453,
    0.04217196, 0.04063930, 0.03910654, 0.03757368, 0.03604074, 0.03450772, 0.03297461, 0.03144142, 0.02990816, 0.02837484,
    0.02684144, 0.02530798, 0.02377446, 0.02224089, 0.02070726, 0.01917358, 0.01763986, 0.01610610, 0.01457230, 0.01303847,
    0.01150460, 0.00997071, 0.00843679, 0.00690286, 0.00536891, 0.00383494, 0.00230097, 0.00076699, -0.00076699, -0.00230097,
    -0.00383494, -0.00536891, -0.00690286, -0.00843679, -0.00997071, -0.01150460, -0.01303847, -0.01457230, -0.01610610, -0.01763986,
    -0.01917358, -0.02070726, -0.02224089, -0.02377446, -0.02530798, -0.02684144, -0.02837484, -0.02990816, -0.03144142, -0.03297461,
    -0.03450772, -0.03604074, -0.03757368, -0.03910654, -0.04063930, -0.04217196, -0.04370453, -0.04523699, -0.04676935, -0.04830159,
    -0.04983373, -0.05136574, -0.05289764, -0.05442941, -0.05596105, -0.05749256, -0.05902393, -0.06055517, -0.06208627, -0.06361721,
    -0.06514801, -0.06667866, -0.06820914, -0.06973947, -0.07126963, -0.07279963, -0.07432945, -0.07585910, -0.07738857, -0.07891786,
    -0.08044697, -0.08197588, -0.08350460, -0.08503312, -0.08656145, -0.08808957, -0.08961748, -0.09114519, -0.09267267, -0.09419994,
    -0.09572699, -0.09725381, -0.09878041, -0.10030677, -0.10183290, -0.10335878, -0.10488442, -0.10640982, -0.10793497, -0.10945986,
    -0.11098449, -0.11250886, -0.11403297, -0.11555681, -0.11708038, -0.11860367, -0.12012669, -0.12164942, -0.12317186, -0.12469402,
    -0.12621588, -0.12773744, -0.12925870, -0.13077966, -0.13230032, -0.13382066, -0.13534068, -0.13686039, -0.13837977, -0.13989883,
    -0.14141756, -0.14293596, -0.14445402, -0.14597174, -0.14748912, -0.14900615, -0.15052283, -0.15203916, -0.15355512, -0.15507073,
    -0.15658597, -0.15810085, -0.15961535, -0.16112947, -0.16264322, -0.16415658, -0.16566956, -0.16718215, -0.16869434, -0.17020614,
    -0.17171754, -0.17322853, -0.17473911, -0.17624929, -0.17775905, -0.17926839, -0.18077731, -0.18228580, -0.18379387, -0.18530150,
    -0.18680870, -0.18831545, -0.18982177, -0.19132763, -0.19283305, -0.19433801, -0.19584252, -0.19734656, -0.19885014, -0.20035326,
    -0.20185590, -0.20335806, -0.20485975, -0.20636096, -0.20786168, -0.20936191, -0.21086164, -0.21236089, -0.21385963, -0.21535787,
    -0.21685560, -0.21835282, -0.21984953, -0.22134572, -0.22284139, -0.22433654, -0.22583115, -0.22732524, -0.22881879, -0.23031180,
    -0.23180428, -0.23329620, -0.23478758, -0.23627840, -0.23776867, -0.23925838, -0.24074752, -0.24223610, -0.24372411, -0.24521155,
    -0.24669841, -0.24818469, -0.24967038, -0.25115549, -0.25264000, -0.25412392, -0.25560725, -0.25708997, -0.25857208, -0.26005359,
    -0.26153449, -0.26301477, -0.26449443, -0.26597347, -0.26745189, -0.26892967, -0.27040682, -0.27188334, -0.27335921, -0.27483445,
    -0.27630903, -0.27778297, -0.27925625, -0.28072887, -0.28220084, -0.28367214, -0.28514277, -0.28661273, -0.28808202, -0.28955063,
    -0.29101856, -0.29248580, -0.29395235, -0.29541822, -0.29688339, -0.29834785, -0.29981162, -0.30127468, -0.30273704, -0.30419868,
    -0.30565960, -0.30711981, -0.30857929, -0.31003805, -0.31149607, -0.31295337, -0.31440993, -0.31586575, -0.31732082, -0.31877515,
    -0.32022873, -0.32168155, -0.32313362, -0.32458492, -0.32603547, -0.32748524, -0.32893425, -0.33038248, -0.33182994, -0.33327661,
    -0.33472250, -0.33616760, -0.33761191, -0.33905543, -0.34049814, -0.34194006, -0.34338117, -0.34482148, -0.34626097, -0.34769965,
    -0.34913751, -0.35057455, -0.35201076, -0.35344614, -0.35488070, -0.35631442, -0.35774730, -0.35917933, -0.36061053, -0.36204087,
    -0.36347036, -0.36489900, -0.36632678, -0.36775370, -0.36917975, -0.37060493, -0.37202924, -0.37345267, -0.37487523, -0.37629691,
    -0.37771769, -0.37913759, -0.38055660, -0.38197471, -0.38339193, -0.38480824, -0.38622364, -0.38763814, -0.38905172, -0.39046439,
    -0.39187614, -0.39328697, -0.39469688, -0.39610585, -0.39751389, -0.39892100, -0.40032717, -0.40173239, -0.40313667, -0.40454000,
    -0.40594238, -0.40734381, -0.40874428, -0.41014378, -0.41154232, -0.41293989, -0.41433649, -0.41573211, -0.41712676, -0.41852043,
    -0.41991310, -0.42130480, -0.42269550, -0.42408520, -0.42547391, -0.42686162, -0.42824832, -0.42963401, -0.43101870, -0.43240237,
    -0.43378502, -0.43516665, -0.43654726, -0.43792683, -0.43930538, -0.44068290, -0.44205938, -0.44343482, -0.44480921, -0.44618256,
    -0.44755486, -0.44892610, -0.45029629, -0.45166542, -0.45303349, -0.45440049, -0.45576642, -0.45713128, -0.45849506, -0.45985776,
    -0.46121939, -0.46257992, -0.46393937, -0.46529773, -0.46665499, -0.46801115, -0.46936622, -0.47072017, -0.47207302, -0.47342476,
    -0.47477539, -0.47612490, -0.47747328, -0.47882055, -0.48016669, -0.48151169, -0.48285557, -0.48419831, -0.48553990, -0.48688036,
    -0.48821967, -0.48955783, -0.49089484, -0.49223070, -0.49356540, -0.49489893, -0.49623130, -0.49756250, -0.49889254, -0.50022139,
    -0.50154908, -0.50287558, -0.50420089, -0.50552503, -0.50684797, -0.50816972, -0.50949027, -0.51080962, -0.51212778, -0.51344472,
    -0.51476046, -0.51607499, -0.51738830, -0.51870040, -0.52001128, -0.52132093, -0.52262935, -0.52393655, -0.52524251, -0.52654724,
    -0.52785072, -0.52915297, -0.53045397, -0.53175372, -0.53305222, -0.53434947, -0.53564546, -0.53694019, -0.53823365, -0.53952585,
    -0.54081678, -0.54210643, -0.54339482, -0.54468192, -0.54596774, -0.54725227, -0.54853552, -0.54981748, -0.55109814, -0.55237751,
    -0.55365558, -0.55493234, -0.55620780, -0.55748195, -0.55875479, -0.56002631, -0.56129651, -0.56256540, -0.56383296, -0.56509919,
    -0.56636410, -0.56762767, -0.56888990, -0.57015080, -0.57141036, -0.57266857, -0.57392543, -0.57518094, -0.57643510, -0.57768790,
    -0.57893935, -0.58018943, -0.58143815, -0.58268549, -0.58393147, -0.58517607, -0.58641930, -0.58766114, -0.58890161, -0.59014068,
    -0.59137837, -0.59261467, -0.59384957, -0.59508308, -0.59631518, -0.59754588, -0.59877518, -0.60000307, -0.60122954, -0.60245460,
    -0.60367824, -0.60490046, -0.60612126, -0.60734063, -0.60855858, -0.60977509, -0.61099016, -0.61220380, -0.61341600, -0.61462676,
    -0.61583606, -0.61704392, -0.61825033, -0.61945528, -0.62065878, -0.62186081, -0.62306138, -0.62426049, -0.62545812, -0.62665429,
    -0.62784898, -0.62904219, -0.63023392, -0.63142417, -0.63261293, -0.63380021, -0.63498599, -0.63617028, -0.63735307, -0.63853436,
    -0.63971415, -0.64089244, -0.64206921, -0.64324448, -0.64441823, -0.64559046, -0.64676118, -0.64793038, -0.64909805, -0.65026419,
    -0.65142880, -0.65259188, -0.65375342, -0.65491343, -0.65607189, -0.65722881, -0.65838419, -0.65953801, -0.66069028, -0.66184100,
    -0.66299016, -0.66413776, -0.66528380, -0.66642827, -0.66757118, -0.66871251, -0.66985227, -0.67099045, -0.67212706, -0.67326208,
    -0.67439552, -0.67552737, -0.67665764, -0.67778631, -0.67891338, -0.68003886, -0.68116274, -0.68228501, -0.68340568, -0.68452474,
    -0.68564219, -0.68675803, -0.68787225, -0.68898485, -0.69009583, -0.69120519, -0.69231292, -0.69341902, -0.69452349, -0.69562633,
    -0.69672753, -0.69782709, -0.69892500, -0.70002128, -0.70111590, -0.70220888, -0.70330020, -0.70438987, -0.70547788, -0.70656423,
    -0.70764892, -0.70873194, -0.70981330, -0.71089298, -0.71197099, -0.71304733, -0.71412199, -0.71519497, -0.71626626, -0.71733587,
    -0.71840380, -0.71947003, -0.72053457, -0.72159741, -0.72265855, -0.72371800, -0.72477574, -0.72583178, -0.72688611, -0.72793872,
    -0.72898963, -0.73003882, -0.73108629, -0.73213204, -0.73317607, -0.73421837, -0.73525895, -0.73629780, -0.73733491, -0.73837029,
    -0.73940393, -0.74043583, -0.74146599, -0.74249440, -0.74352107, -0.74454598, -0.74556915, -0.74659056, -0.74761021, -0.74862811,
    -0.74964424, -0.75065861, -0.75167121, -0.75268205, -0.75369111, -0.75469840, -0.75570391, -0.75670765, -0.75770960, -0.75870977,
    -0.75970816, -0.76070476, -0.76169957, -0.76269258, -0.76368380, -0.76467323, -0.76566085, -0.76664668, -0.76763070, -0.76861291,
    -0.76959331, -0.77057191, -0.77154869, -0.77252365, -0.77349680, -0.77446813, -0.77543763, -0.77640531, -0.77737116, -0.77833519,
    -0.77929738, -0.78025774, -0.78121626, -0.78217294, -0.78312779, -0.78408079, -0.78503194, -0.78598125, -0.78692871, -0.78787432,
    -0.78881807, -0.78975997, -0.79070001, -0.79163819, -0.79257450, -0.79350895, -0.79444154, -0.79537225, -0.79630109, -0.79722806,
    -0.79815315, -0.79907637, -0.79999770, -0.80091715, -0.80183472, -0.80275040, -0.80366419, -0.80457609, -0.80548610, -0.80639421,
    -0.80730042, -0.80820474, -0.80910715, -0.81000766, -0.81090626, -0.81180296, -0.81269774, -0.81359061, -0.81448157, -0.81537061,
    -0.81625773, -0.81714293, -0.81802621, -0.81890757, -0.81978699, -0.82066449, -0.82154006, -0.82241369, -0.82328539, -0.82415515,
    -0.82502297, -0.82588885, -0.82675279, -0.82761478, -0.82847482, -0.82933292, -0.83018906, -0.83104325, -0.83189548, -0.83274576,
    -0.83359408, -0.83444043, -0.83528483, -0.83612725, -0.83696771, -0.83780620, -0.83864272, -0.83947726, -0.84030983, -0.84114042,
    -0.84196904, -0.84279567, -0.84362032, -0.84444298, -0.84526365, -0.84608234, -0.84689904, -0.84771374, -0.84852645, -0.84933716,
    -0.85014587, -0.85095259, -0.85175730, -0.85256000, -0.85336070, -0.85415940, -0.85495608, -0.85575075, -0.85654340, -0.85733405,
    -0.85812267, -0.85890927, -0.85969386, -0.86047642, -0.86125695, -0.86203546, -0.86281194, -0.86358639, -0.86435881, -0.86512920,
    -0.86589754, -0.86666385, -0.86742813, -0.86819036, -0.86895054, -0.86970869, -0.87046478, -0.87121883, -0.87197083, -0.87272078,
    -0.87346867, -0.87421451, -0.87495829, -0.87570001, -0.87643967, -0.87717727, -0.87791280, -0.87864627, -0.87937767, -0.88010700,
    -0.88083426, -0.88155945, -0.88228256, -0.88300360, -0.88372256, -0.88443944, -0.88515424, -0.88586695, -0.88657759, -0.88728613,
    -0.88799259, -0.88869696, -0.88939923, -0.89009942, -0.89079751, -0.89149350, -0.89218739, -0.89287919, -0.89356889, -0.89425648,
    -0.89494197, -0.89562535, -0.89630662, -0.89698579, -0.89766284, -0.89833779, -0.89901062, -0.89968133, -0.90034993, -0.90101640,
    -0.90168076, -0.90234300, -0.90300311, -0.90366110, -0.90431696, -0.90497069, -0.90562229, -0.90627177, -0.90691911, -0.90756431,
    -0.90820738, -0.90884832, -0.90948711, -0.91012377, -0.91075828, -0.91139065, -0.91202088, -0.91264896, -0.91327489, -0.91389867,
    -0.91452030, -0.91513978, -0.91575711, -0.91637228, -0.91698530, -0.91759616, -0.91820486, -0.91881139, -0.91941577, -0.92001798,
    -0.92061803, -0.92121591, -0.92181163, -0.92240517, -0.92299654, -0.92358575, -0.92417278, -0.92475763, -0.92534031, -0.92592081,
    -0.92649913, -0.92707527, -0.92764923, -0.92822101, -0.92879060, -0.92935801, -0.92992323, -0.93048627, -0.93104711, -0.93160576,
    -0.93216222, -0.93271649, -0.93326856, -0.93381844, -0.93436611, -0.93491159, -0.93545487, -0.93599595, -0.93653483, -0.93707150,
    -0.93760597, -0.93813823, -0.93866828, -0.93919613, -0.93972176, -0.94024519, -0.94076640, -0.94128540, -0.94180218, -0.94231675,
    -0.94282909, -0.94333923, -0.94384714, -0.94435283, -0.94485629, -0.94535754, -0.94585656, -0.94635335, -0.94684792, -0.94734026,
    -0.94783037, -0.94831825, -0.94880389, -0.94928731, -0.94976849, -0.95024744, -0.95072415, -0.95119862, -0.95167086, -0.95214085,
    -0.95260861, -0.95307412, -0.95353740, -0.95399842, -0.95445721, -0.95491374, -0.95536803, -0.95582007, -0.95626987, -0.95671741,
    -0.95716270, -0.95760574, -0.95804652, -0.95848506, -0.95892133, -0.95935535, -0.95978711, -0.96021662, -0.96064386, -0.96106884,
    -0.96149156, -0.96191202, -0.96233022, -0.96274615, -0.96315982, -0.96357122, -0.96398035, -0.96438721, -0.96479181, -0.96519413,
    -0.96559418, -0.96599197, -0.96638747, -0.96678071, -0.96717167, -0.96756035, -0.96794676, -0.96833088, -0.96871273, -0.96909231,
    -0.96946960, -0.96984460, -0.97021733, -0.97058778, -0.97095594, -0.97132181, -0.97168540, -0.97204670, -0.97240572, -0.97276245,
    -0.97311689, -0.97346903, -0.97381889, -0.97416646, -0.97451173, -0.97485471, -0.97519540, -0.97553379, -0.97586989, -0.97620369,
    -0.97653520, -0.97686440, -0.97719131, -0.97751592, -0.97783822, -0.97815823, -0.97847594, -0.97879134, -0.97910444, -0.97941523,
    -0.97972372, -0.98002991, -0.98033379, -0.98063536, -0.98093462, -0.98123158, -0.98152623, -0.98181857, -0.98210859, -0.98239631,
    -0.98268172, -0.98296481, -0.98324559, -0.98352405, -0.98380021, -0.98407404, -0.98434556, -0.98461477, -0.98488166, -0.98514623,
    -0.98540848, -0.98566841, -0.98592603, -0.98618132, -0.98643429, -0.98668495, -0.98693328, -0.98717929, -0.98742297, -0.98766433,
    -0.98790337, -0.98814008, -0.98837447, -0.98860653, -0.98883627, -0.98906368, -0.98928876, -0.98951151, -0.98973194, -0.98995004,
    -0.99016580, -0.99037924, -0.99059035, -0.99079912, -0.99100557, -0.99120968, -0.99141146, -0.99161091, -0.99180802, -0.99200280,
    -0.99219524, -0.99238535, -0.99257313, -0.99275857, -0.99294167, -0.99312244, -0.99330087, -0.99347697, -0.99365072, -0.99382214,
    -0.99399122, -0.99415796, -0.99432236, -0.99448442, -0.99464414, -0.99480152, -0.99495656, -0.99510926, -0.99525961, -0.99540763,
    -0.99555330, -0.99569663, -0.99583761, -0.99597626, -0.99611256, -0.99624651, -0.99637812, -0.99650739, -0.99663431, -0.99675889,
    -0.99688112, -0.99700101, -0.99711855, -0.99723374, -0.99734659, -0.99745709, -0.99756524, -0.99767104, -0.99777450, -0.99787561,
    -0.99797437, -0.99807079, -0.99816485, -0.99825657, -0.99834593, -0.99843295, -0.99851762, -0.99859994, -0.99867991, -0.99875753,
    -0.99883280, -0.99890572, -0.99897628, -0.99904450, -0.99911037, -0.99917388, -0.99923505, -0.99929386, -0.99935032, -0.99940443,
    -0.99945619, -0.99950560, -0.99955265, -0.99959735, -0.99963970, -0.99967970, -0.99971735, -0.99975264, -0.99978558, -0.99981617,
    -0.99984441, -0.99987029, -0.99989382, -0.99991500, -0.99993382, -0.99995029, -0.99996441, -0.99997617, -0.99998559, -0.99999265,
    -0.99999735, -0.99999971, -0.99999971, -0.99999735, -0.99999265, -0.99998559, -0.99997617, -0.99996441, -0.99995029, -0.99993382,
    -0.99991500, -0.99989382, -0.99987029, -0.99984441, -0.99981617, -0.99978558, -0.99975264, -0.99971735, -0.99967970, -0.99963970,
    -0.99959735, -0.99955265, -0.99950560, -0.99945619, -0.99940443, -0.99935032, -0.99929386, -0.99923505, -0.99917388, -0.99911037,
    -0.99904450, -0.99897628, -0.99890572, -0.99883280, -0.99875753, -0.99867991, -0.99859994, -0.99851762, -0.99843295, -0.99834593,
    -0.99825657, -0.99816485, -0.99807079, -0.99797437, -0.99787561, -0.99777450, -0.99767104, -0.99756524, -0.99745709, -0.99734659,
    -0.99723374, -0.99711855, -0.99700101, -0.99688112, -0.99675889, -0.99663431, -0.99650739, -0.99637812, -0.99624651, -0.99611256,
    -0.99597626, -0.99583761, -0.99569663, -0.99555330, -0.99540763, -0.99525961, -0.99510926, -0.99495656, -0.99480152, -0.99464414,
    -0.99448442, -0.99432236, -0.99415796, -0.99399122, -0.99382214, -0.99365072, -0.99347697, -0.99330087, -0.99312244, -0.99294167,
    -0.99275857, -0.99257313, -0.99238535, -0.99219524, -0.99200280, -0.99180802, -0.99161091, -0.99141146, -0.99120968, -0.99100557,
    -0.99079912, -0.99059035, -0.99037924, -0.99016580, -0.98995004, -0.98973194, -0.98951151, -0.98928876, -0.98906368, -0.98883627,
    -0.98860653, -0.98837447, -0.98814008, -0.98790337, -0.98766433, -0.98742297, -0.98717929, -0.98693328, -0.98668495, -0.98643429,
    -0.98618132, -0.98592603, -0.98566841, -0.98540848, -0.98514623, -0.98488166, -0.98461477, -0.98434556, -0.98407404, -0.98380021,
    -0.98352405, -0.98324559, -0.98296481, -0.98268172, -0.98239631, -0.98210859, -0.98181857, -0.98152623, -0.98123158, -0.98093462,
    -0.98063536, -0.98033379, -0.98002991, -0.97972372, -0.97941523, -0.97910444, -0.97879134, -0.97847594, -0.97815823, -0.97783822,
    -0.97751592, -0.97719131, -0.97686440, -0.97653520, -0.97620369, -0.97586989, -0.97553379, -0.97519540, -0.97485471, -0.97451173,
    -0.97416646, -0.97381889, -0.97346903, -0.97311689, -0.97276245, -0.97240572, -0.97204670, -0.97168540, -0.97132181, -0.97095594,
    -0.97058778, -0.97021733, -0.96984460, -0.96946960, -0.96909231, -0.96871273, -0.96833088, -0.96794676, -0.96756035, -0.96717167,
    -0.96678071, -0.96638747, -0.96599197, -0.96559418, -0.96519413, -0.96479181, -0.96438721, -0.96398035, -0.96357122, -0.96315982,
    -0.96274615, -0.96233022, -0.96191202, -0.96149156, -0.96106884, -0.96064386, -0.96021662, -0.95978711, -0.95935535, -0.95892133,
    -0.95848506, -0.95804652, -0.95760574, -0.95716270, -0.95671741, -0.95626987, -0.95582007, -0.95536803, -0.95491374, -0.95445721,
    -0.95399842, -0.95353740, -0.95307412, -0.95260861, -0.95214085, -0.95167086, -0.95119862, -0.95072415, -0.95024744, -0.94976849,
    -0.94928731, -0.94880389, -0.94831825, -0.94783037, -0.94734026, -0.94684792, -0.94635335, -0.94585656, -0.94535754, -0.94485629,
    -0.94435283, -0.94384714, -0.94333923, -0.94282909, -0.94231675, -0.94180218, -0.94128540, -0.94076640, -0.94024519, -0.93972176,
    -0.93919613, -0.93866828, -0.93813823, -0.93760597, -0.93707150, -0.93653483, -0.93599595, -0.93545487, -0.93491159, -0.93436611,
    -0.93381844, -0.93326856, -0.93271649, -0.93216222, -0.93160576, -0.93104711, -0.93048627, -0.92992323, -0.92935801, -0.92879060,
    -0.92822101, -0.92764923, -0.92707527, -0.92649913, -0.92592081, -0.92534031, -0.92475763, -0.92417278, -0.92358575, -0.92299654,
    -0.92240517, -0.92181163, -0.92121591, -0.92061803, -0.92001798, -0.91941577, -0.91881139, -0.91820486, -0.91759616, -0.91698530,
    -0.91637228, -0.91575711, -0.91513978, -0.91452030, -0.91389867, -0.91327489, -0.91264896, -0.91202088, -0.91139065, -0.91075828,
    -0.91012377, -0.90948711, -0.90884832, -0.90820738, -0.90756431, -0.90691911, -0.90627177, -0.90562229, -0.90497069, -0.90431696,
    -0.90366110, -0.90300311, -0.90234300, -0.90168076, -0.90101640, -0.90034993, -0.89968133, -0.89901062, -0.89833779, -0.89766284,
    -0.89698579, -0.89630662, -0.89562535, -0.89494197, -0.89425648, -0.89356889, -0.89287919, -0.89218739, -0.89149350, -0.89079751,
    -0.89009942, -0.88939923, -0.88869696, -0.88799259, -0.88728613, -0.88657759, -0.88586695, -0.88515424, -0.88443944, -0.88372256,
    -0.88300360, -0.88228256, -0.88155945, -0.88083426, -0.88010700, -0.87937767, -0.87864627, -0.87791280, -0.87717727, -0.87643967,
    -0.87570001, -0.87495829, -0.87421451, -0.87346867, -0.87272078, -0.87197083, -0.87121883, -0.87046478, -0.86970869, -0.86895054,
    -0.86819036, -0.86742813, -0.86666385, -0.86589754, -0.86512920, -0.86435881, -0.86358639, -0.86281194, -0.86203546, -0.86125695,
    -0.86047642, -0.85969386, -0.85890927, -0.85812267, -0.85733405, -0.85654340, -0.85575075, -0.85495608, -0.85415940, -0.85336070,
    -0.85256000, -0.85175730, -0.85095259, -0.85014587, -0.84933716, -0.84852645, -0.84771374, -0.84689904, -0.84608234, -0.84526365,
    -0.84444298, -0.84362032, -0.84279567, -0.84196904, -0.84114042, -0.84030983, -0.83947726, -0.83864272, -0.83780620, -0.83696771,
    -0.83612725, -0.83528483, -0.83444043, -0.83359408, -0.83274576, -0.83189548, -0.83104325, -0.83018906, -0.82933292, -0.82847482,
    -0.82761478, -0.82675279, -0.82588885, -0.82502297, -0.82415515, -0.82328539, -0.82241369, -0.82154006, -0.82066449, -0.81978699,
    -0.81890757, -0.81802621, -0.81714293, -0.81625773, -0.81537061, -0.81448157, -0.81359061, -0.81269774, -0.81180296, -0.81090626,
    -0.81000766, -0.80910715, -0.80820474, -0.80730042, -0.80639421, -0.80548610, -0.80457609, -0.80366419, -0.80275040, -0.80183472,
    -0.80091715, -0.79999770, -0.79907637, -0.79815315, -0.79722806, -0.79630109, -0.79537225, -0.79444154, -0.79350895, -0.79257450,
    -0.79163819, -0.79070001, -0.78975997, -0.78881807, -0.78787432, -0.78692871, -0.78598125, -0.78503194, -0.78408079, -0.78312779,
    -0.78217294, -0.78121626, -0.78025774, -0.77929738, -0.77833519, -0.77737116, -0.77640531, -0.77543763, -0.77446813, -0.77349680,
    -0.77252365, -0.77154869, -0.77057191, -0.76959331, -0.76861291, -0.76763070, -0.76664668, -0.76566085, -0.76467323, -0.76368380,
    -0.76269258, -0.76169957, -0.76070476, -0.75970816, -0.75870977, -0.75770960, -0.75670765, -0.75570391, -0.75469840, -0.75369111,
    -0.75268205, -0.75167121, -0.75065861, -0.74964424, -0.74862811, -0.74761021, -0.74659056, -0.74556915, -0.74454598, -0.74352107,
    -0.74249440, -0.74146599, -0.74043583, -0.73940393, -0.73837029, -0.73733491, -0.73629780, -0.73525895, -0.73421837, -0.73317607,
    -0.73213204, -0.73108629, -0.73003882, -0.72898963, -0.72793872, -0.72688611, -0.72583178, -0.72477574, -0.72371800, -0.72265855,
    -0.72159741, -0.72053457, -0.71947003, -0.71840380, -0.71733587, -0.71626626, -0.71519497, -0.71412199, -0.71304733, -0.71197099,
    -0.71089298, -0.70981330, -0.70873194, -0.70764892, -0.70656423, -0.70547788, -0.70438987, -0.70330020, -0.70220888, -0.70111590,
    -0.70002128, -0.69892500, -0.69782709, -0.69672753, -0.69562633, -0.69452349, -0.69341902, -0.69231292, -0.69120519, -0.69009583,
    -0.68898485, -0.68787225, -0.68675803, -0.68564219, -0.68452474, -0.68340568, -0.68228501, -0.68116274, -0.68003886, -0.67891338,
    -0.67778631, -0.67665764, -0.67552737, -0.67439552, -0.67326208, -0.67212706, -0.67099045, -0.66985227, -0.66871251, -0.66757118,
    -0.66642827, -0.66528380, -0.66413776, -0.66299016, -0.66184100, -0.66069028, -0.65953801, -0.65838419, -0.65722881, -0.65607189,
    -0.65491343, -0.65375342, -0.65259188, -0.65142880, -0.65026419, -0.64909805, -0.64793038, -0.64676118, -0.64559046, -0.64441823,
    -0.64324448, -0.64206921, -0.64089244, -0.63971415, -0.63853436, -0.63735307, -0.63617028, -0.63498599, -0.63380021, -0.63261293,
    -0.63142417, -0.63023392, -0.62904219, -0.62784898, -0.62665429, -0.62545812, -0.62426049, -0.62306138, -0.62186081, -0.62065878,
    -0.61945528, -0.61825033, -0.61704392, -0.61583606, -0.61462676, -0.61341600, -0.61220380, -0.61099016, -0.60977509, -0.60855858,
    -0.60734063, -0.60612126, -0.60490046, -0.60367824, -0.60245460, -0.60122954, -0.60000307, -0.59877518, -0.59754588, -0.59631518,
    -0.59508308, -0.59384957, -0.59261467, -0.59137837, -0.59014068, -0.58890161, -0.58766114, -0.58641930, -0.58517607, -0.58393147,
    -0.58268549, -0.58143815, -0.58018943, -0.57893935, -0.57768790, -0.57643510, -0.57518094, -0.57392543, -0.57266857, -0.57141036,
    -0.57015080, -0.56888990, -0.56762767, -0.56636410, -0.56509919, -0.56383296, -0.56256540, -0.56129651, -0.56002631, -0.55875479,
    -0.55748195, -0.55620780, -0.55493234, -0.55365558, -0.55237751, -0.55109814, -0.54981748, -0.54853552, -0.54725227, -0.54596774,
    -0.54468192, -0.54339482, -0.54210643, -0.54081678, -0.53952585, -0.53823365, -0.53694019, -0.53564546, -0.53434947, -0.53305222,
    -0.53175372, -0.53045397, -0.52915297, -0.52785072, -0.52654724, -0.52524251, -0.52393655, -0.52262935, -0.52132093, -0.52001128,
    -0.51870040, -0.51738830, -0.51607499, -0.51476046, -0.51344472, -0.51212778, -0.51080962, -0.50949027, -0.50816972, -0.50684797,
    -0.50552503, -0.50420089, -0.50287558, -0.50154908, -0.50022139, -0.49889254, -0.49756250, -0.49623130, -0.49489893, -0.49356540,
    -0.49223070, -0.49089484, -0.48955783, -0.48821967, -0.48688036, -0.48553990, -0.48419831, -0.48285557, -0.48151169, -0.48016669,
    -0.47882055, -0.47747328, -0.47612490, -0.47477539, -0.47342476, -0.47207302, -0.47072017, -0.46936622, -0.46801115, -0.46665499,
    -0.46529773, -0.46393937, -0.46257992, -0.46121939, -0.45985776, -0.45849506, -0.45713128, -0.45576642, -0.45440049, -0.45303349,
    -0.45166542, -0.45029629, -0.44892610, -0.44755486, -0.44618256, -0.44480921, -0.44343482, -0.44205938, -0.44068290, -0.43930538,
    -0.43792683, -0.43654726, -0.43516665, -0.43378502, -0.43240237, -0.43101870, -0.42963401, -0.42824832, -0.42686162, -0.42547391,
    -0.42408520, -0.42269550, -0.42130480, -0.41991310, -0.41852043, -0.41712676, -0.41573211, -0.41433649, -0.41293989, -0.41154232,
    -0.41014378, -0.40874428, -0.40734381, -0.40594238, -0.40454000, -0.40313667, -0.40173239, -0.40032717, -0.39892100, -0.39751389,
    -0.39610585, -0.39469688, -0.39328697, -0.39187614, -0.39046439, -0.38905172, -0.38763814, -0.38622364, -0.38480824, -0.38339193,
    -0.38197471, -0.38055660, -0.37913759, -0.37771769, -0.37629691, -0.37487523, -0.37345267, -0.37202924, -0.37060493, -0.36917975,
    -0.36775370, -0.36632678, -0.36489900, -0.36347036, -0.36204087, -0.36061053, -0.35917933, -0.35774730, -0.35631442, -0.35488070,
    -0.35344614, -0.35201076, -0.35057455, -0.34913751, -0.34769965, -0.34626097, -0.34482148, -0.34338117, -0.34194006, -0.34049814,
    -0.33905543, -0.33761191, -0.33616760, -0.33472250, -0.33327661, -0.33182994, -0.33038248, -0.32893425, -0.32748524, -0.32603547,
    -0.32458492, -0.32313362, -0.32168155, -0.32022873, -0.31877515, -0.31732082, -0.31586575, -0.31440993, -0.31295337, -0.31149607,
    -0.31003805, -0.30857929, -0.30711981, -0.30565960, -0.30419868, -0.30273704, -0.30127468, -0.29981162, -0.29834785, -0.29688339,
    -0.29541822, -0.29395235, -0.29248580, -0.29101856, -0.28955063, -0.28808202, -0.28661273, -0.28514277, -0.28367214, -0.28220084,
    -0.28072887, -0.27925625, -0.27778297, -0.27630903, -0.27483445, -0.27335921, -0.27188334, -0.27040682, -0.26892967, -0.26745189,
    -0.26597347, -0.26449443, -0.26301477, -0.26153449, -0.26005359, -0.25857208, -0.25708997, -0.25560725, -0.25412392, -0.25264000,
    -0.25115549, -0.24967038, -0.24818469, -0.24669841, -0.24521155, -0.24372411, -0.24223610, -0.24074752, -0.23925838, -0.23776867,
    -0.23627840, -0.23478758, -0.23329620, -0.23180428, -0.23031180, -0.22881879, -0.22732524, -0.22583115, -0.22433654, -0.22284139,
    -0.22134572, -0.21984953, -0.21835282, -0.21685560, -0.21535787, -0.21385963, -0.21236089, -0.21086164, -0.20936191, -0.20786168,
    -0.20636096, -0.20485975, -0.20335806, -0.20185590, -0.20035326, -0.19885014, -0.19734656, -0.19584252, -0.19433801, -0.19283305,
    -0.19132763, -0.18982177, -0.18831545, -0.18680870, -0.18530150, -0.18379387, -0.18228580, -0.18077731, -0.17926839, -0.17775905,
    -0.17624929, -0.17473911, -0.17322853, -0.17171754, -0.17020614, -0.16869434, -0.16718215, -0.16566956, -0.16415658, -0.16264322,
    -0.16112947, -0.15961535, -0.15810085, -0.15658597, -0.15507073, -0.15355512, -0.15203916, -0.15052283, -0.14900615, -0.14748912,
    -0.14597174, -0.14445402, -0.14293596, -0.14141756, -0.13989883, -0.13837977, -0.13686039, -0.13534068, -0.13382066, -0.13230032,
    -0.13077966, -0.12925870, -0.12773744, -0.12621588, -0.12469402, -0.12317186, -0.12164942, -0.12012669, -0.11860367, -0.11708038,
    -0.11555681, -0.11403297, -0.11250886, -0.11098449, -0.10945986, -0.10793497, -0.10640982, -0.10488442, -0.10335878, -0.10183290,
    -0.10030677, -0.09878041, -0.09725381, -0.09572699, -0.09419994, -0.09267267, -0.09114519, -0.08961748, -0.08808957, -0.08656145,
    -0.08503312, -0.08350460, -0.08197588, -0.08044697, -0.07891786, -0.07738857, -0.07585910, -0.07432945, -0.07279963, -0.07126963,
    -0.06973947, -0.06820914, -0.06667866, -0.06514801, -0.06361721, -0.06208627, -0.06055517, -0.05902393, -0.05749256, -0.05596105,
    -0.05442941, -0.05289764, -0.05136574, -0.04983373, -0.04830159, -0.04676935, -0.04523699, -0.04370453, -0.04217196, -0.04063930,
    -0.03910654, -0.03757368, -0.03604074, -0.03450772, -0.03297461, -0.03144142, -0.02990816, -0.02837484, -0.02684144, -0.02530798,
    -0.02377446, -0.02224089, -0.02070726, -0.01917358, -0.01763986, -0.01610610, -0.01457230, -0.01303847, -0.01150460, -0.00997071,
    -0.00843679, -0.00690286, -0.00536891, -0.00383494, -0.00230097, -0.00076699
    );

end package sin_4096;
