-------------------------------------------------------------------------------
-- Title       : Testbench Equalizer
-- Author      : Michael Wurm <michael.wurm@students.fh-hagenberg.at>
-------------------------------------------------------------------------------
-- Description : Bandpasses equally distributed on frequency range (10Hz-20kHz)
--               each with a configurable factor
-------------------------------------------------------------------------------

entity tbEqualizer is
end entity tbEqualizer;

architecture bhv of tbEqualizer is
    ---------------------------------------------------------------------------
    -- Constants
    ---------------------------------------------------------------------------

    ---------------------------------------------------------------------------
    -- Signals
    ---------------------------------------------------------------------------

begin

    ---------------------------------------------------------------------------
    -- Signal assignments
    ---------------------------------------------------------------------------
    Clk <= not Clk after 10 ns;

    ---------------------------------------------------------------------------
    -- Instantiations
    ---------------------------------------------------------------------------

end architecture bhv;
