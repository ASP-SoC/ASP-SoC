architecture Struct of AudioCodecAvalon is

begin  -- architecture Struct

  

end architecture Struct;
