-- Audio.vhd

-- Generated using ACDS version 16.1 203

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Audio is
	port (
		audio_clk_clk : out   std_logic;        -- audio_clk.clk
		clk_clk       : in    std_logic := '0'; --       clk.clk
		i2c_SDAT      : inout std_logic := '0'; --       i2c.SDAT
		i2c_SCLK      : out   std_logic;        --          .SCLK
		i2s_adcdat    : in    std_logic := '0'; --       i2s.adcdat
		i2s_adclrck   : in    std_logic := '0'; --          .adclrck
		i2s_bclk      : in    std_logic := '0'; --          .bclk
		i2s_dacdat    : out   std_logic;        --          .dacdat
		i2s_daclrck   : in    std_logic := '0'; --          .daclrck
		reset_reset_n : in    std_logic := '0'  --     reset.reset_n
	);
end entity Audio;

architecture rtl of Audio is
	component AudioCodecAvalon is
		generic (
			gDataWidth    : natural := 24;
			gDataWidthLen : natural := 5
		);
		port (
			csi_clk         : in  std_logic                     := 'X';             -- clk
			rsi_reset_n     : in  std_logic                     := 'X';             -- reset_n
			AUD_ADCDAT      : in  std_logic                     := 'X';             -- adcdat
			AUD_ADCLRCK     : in  std_logic                     := 'X';             -- adclrck
			AUD_BCLK        : in  std_logic                     := 'X';             -- bclk
			AUD_DACDAT      : out std_logic;                                        -- dacdat
			AUD_DACLRCK     : in  std_logic                     := 'X';             -- daclrck
			asi_left_data   : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			asi_left_valid  : in  std_logic                     := 'X';             -- valid
			asi_right_data  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			asi_right_valid : in  std_logic                     := 'X';             -- valid
			aso_left_data   : out std_logic_vector(23 downto 0);                    -- data
			aso_left_valid  : out std_logic;                                        -- valid
			aso_right_data  : out std_logic_vector(23 downto 0);                    -- data
			aso_right_valid : out std_logic                                         -- valid
		);
	end component AudioCodecAvalon;

	component FIR is
		generic (
			gDataWidth      : natural := 24;
			gNrAddressLines : natural := 4
		);
		port (
			csi_clk          : in  std_logic                     := 'X';             -- clk
			rsi_reset_n      : in  std_logic                     := 'X';             -- reset_n
			avs_s0_address   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			avs_s0_write     : in  std_logic                     := 'X';             -- write
			avs_s0_writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_s0_read      : in  std_logic                     := 'X';             -- read
			avs_s0_readdata  : out std_logic_vector(31 downto 0);                    -- readdata
			asi_valid        : in  std_logic                     := 'X';             -- valid
			asi_data         : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			aso_valid        : out std_logic;                                        -- valid
			aso_data         : out std_logic_vector(23 downto 0)                     -- data
		);
	end component FIR;

	component Audio_audio_config is
		port (
			clk         : in    std_logic                     := 'X';             -- clk
			reset       : in    std_logic                     := 'X';             -- reset
			address     : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable  : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			read        : in    std_logic                     := 'X';             -- read
			write       : in    std_logic                     := 'X';             -- write
			writedata   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata    : out   std_logic_vector(31 downto 0);                    -- readdata
			waitrequest : out   std_logic;                                        -- waitrequest
			I2C_SDAT    : inout std_logic                     := 'X';             -- export
			I2C_SCLK    : out   std_logic                                         -- export
		);
	end component Audio_audio_config;

	component Audio_audio_pll is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			audio_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component Audio_audio_pll;

	component Audio_jtag is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component Audio_jtag;

	component Audio_nios is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(13 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(13 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component Audio_nios;

	component Audio_onchip_memory is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component Audio_onchip_memory;

	component Audio_mm_interconnect_0 is
		port (
			clk_clk_clk                            : in  std_logic                     := 'X';             -- clk
			nios_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios_data_master_address               : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			nios_data_master_waitrequest           : out std_logic;                                        -- waitrequest
			nios_data_master_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios_data_master_read                  : in  std_logic                     := 'X';             -- read
			nios_data_master_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			nios_data_master_write                 : in  std_logic                     := 'X';             -- write
			nios_data_master_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios_data_master_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			nios_instruction_master_address        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			nios_instruction_master_waitrequest    : out std_logic;                                        -- waitrequest
			nios_instruction_master_read           : in  std_logic                     := 'X';             -- read
			nios_instruction_master_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			Avalon_FIR_0_s0_address                : out std_logic_vector(3 downto 0);                     -- address
			Avalon_FIR_0_s0_write                  : out std_logic;                                        -- write
			Avalon_FIR_0_s0_read                   : out std_logic;                                        -- read
			Avalon_FIR_0_s0_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Avalon_FIR_0_s0_writedata              : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_avalon_jtag_slave_address         : out std_logic_vector(0 downto 0);                     -- address
			jtag_avalon_jtag_slave_write           : out std_logic;                                        -- write
			jtag_avalon_jtag_slave_read            : out std_logic;                                        -- read
			jtag_avalon_jtag_slave_readdata        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_avalon_jtag_slave_writedata       : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_avalon_jtag_slave_waitrequest     : in  std_logic                     := 'X';             -- waitrequest
			jtag_avalon_jtag_slave_chipselect      : out std_logic;                                        -- chipselect
			nios_debug_mem_slave_address           : out std_logic_vector(8 downto 0);                     -- address
			nios_debug_mem_slave_write             : out std_logic;                                        -- write
			nios_debug_mem_slave_read              : out std_logic;                                        -- read
			nios_debug_mem_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios_debug_mem_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			nios_debug_mem_slave_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			nios_debug_mem_slave_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			nios_debug_mem_slave_debugaccess       : out std_logic;                                        -- debugaccess
			onchip_memory_s1_address               : out std_logic_vector(9 downto 0);                     -- address
			onchip_memory_s1_write                 : out std_logic;                                        -- write
			onchip_memory_s1_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory_s1_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory_s1_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory_s1_chipselect            : out std_logic;                                        -- chipselect
			onchip_memory_s1_clken                 : out std_logic                                         -- clken
		);
	end component Audio_mm_interconnect_0;

	component Audio_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component Audio_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal avalon_fir_0_avalon_streaming_source_0_valid             : std_logic;                     -- Avalon_FIR_0:aso_valid -> AudioCodecAvalon_0:asi_left_valid
	signal avalon_fir_0_avalon_streaming_source_0_data              : std_logic_vector(23 downto 0); -- Avalon_FIR_0:aso_data -> AudioCodecAvalon_0:asi_left_data
	signal audiocodecavalon_0_left_source_valid                     : std_logic;                     -- AudioCodecAvalon_0:aso_left_valid -> Avalon_FIR_0:asi_valid
	signal audiocodecavalon_0_left_source_data                      : std_logic_vector(23 downto 0); -- AudioCodecAvalon_0:aso_left_data -> Avalon_FIR_0:asi_data
	signal audiocodecavalon_0_right_source_valid                    : std_logic;                     -- AudioCodecAvalon_0:aso_right_valid -> AudioCodecAvalon_0:asi_right_valid
	signal audiocodecavalon_0_right_source_data                     : std_logic_vector(23 downto 0); -- AudioCodecAvalon_0:aso_right_data -> AudioCodecAvalon_0:asi_right_data
	signal nios_data_master_readdata                                : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios_data_master_readdata -> nios:d_readdata
	signal nios_data_master_waitrequest                             : std_logic;                     -- mm_interconnect_0:nios_data_master_waitrequest -> nios:d_waitrequest
	signal nios_data_master_debugaccess                             : std_logic;                     -- nios:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios_data_master_debugaccess
	signal nios_data_master_address                                 : std_logic_vector(13 downto 0); -- nios:d_address -> mm_interconnect_0:nios_data_master_address
	signal nios_data_master_byteenable                              : std_logic_vector(3 downto 0);  -- nios:d_byteenable -> mm_interconnect_0:nios_data_master_byteenable
	signal nios_data_master_read                                    : std_logic;                     -- nios:d_read -> mm_interconnect_0:nios_data_master_read
	signal nios_data_master_write                                   : std_logic;                     -- nios:d_write -> mm_interconnect_0:nios_data_master_write
	signal nios_data_master_writedata                               : std_logic_vector(31 downto 0); -- nios:d_writedata -> mm_interconnect_0:nios_data_master_writedata
	signal nios_instruction_master_readdata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios_instruction_master_readdata -> nios:i_readdata
	signal nios_instruction_master_waitrequest                      : std_logic;                     -- mm_interconnect_0:nios_instruction_master_waitrequest -> nios:i_waitrequest
	signal nios_instruction_master_address                          : std_logic_vector(13 downto 0); -- nios:i_address -> mm_interconnect_0:nios_instruction_master_address
	signal nios_instruction_master_read                             : std_logic;                     -- nios:i_read -> mm_interconnect_0:nios_instruction_master_read
	signal mm_interconnect_0_nios_debug_mem_slave_readdata          : std_logic_vector(31 downto 0); -- nios:debug_mem_slave_readdata -> mm_interconnect_0:nios_debug_mem_slave_readdata
	signal mm_interconnect_0_nios_debug_mem_slave_waitrequest       : std_logic;                     -- nios:debug_mem_slave_waitrequest -> mm_interconnect_0:nios_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios_debug_mem_slave_debugaccess       : std_logic;                     -- mm_interconnect_0:nios_debug_mem_slave_debugaccess -> nios:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios_debug_mem_slave_address           : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios_debug_mem_slave_address -> nios:debug_mem_slave_address
	signal mm_interconnect_0_nios_debug_mem_slave_read              : std_logic;                     -- mm_interconnect_0:nios_debug_mem_slave_read -> nios:debug_mem_slave_read
	signal mm_interconnect_0_nios_debug_mem_slave_byteenable        : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios_debug_mem_slave_byteenable -> nios:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios_debug_mem_slave_write             : std_logic;                     -- mm_interconnect_0:nios_debug_mem_slave_write -> nios:debug_mem_slave_write
	signal mm_interconnect_0_nios_debug_mem_slave_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios_debug_mem_slave_writedata -> nios:debug_mem_slave_writedata
	signal mm_interconnect_0_avalon_fir_0_s0_readdata               : std_logic_vector(31 downto 0); -- Avalon_FIR_0:avs_s0_readdata -> mm_interconnect_0:Avalon_FIR_0_s0_readdata
	signal mm_interconnect_0_avalon_fir_0_s0_address                : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Avalon_FIR_0_s0_address -> Avalon_FIR_0:avs_s0_address
	signal mm_interconnect_0_avalon_fir_0_s0_read                   : std_logic;                     -- mm_interconnect_0:Avalon_FIR_0_s0_read -> Avalon_FIR_0:avs_s0_read
	signal mm_interconnect_0_avalon_fir_0_s0_write                  : std_logic;                     -- mm_interconnect_0:Avalon_FIR_0_s0_write -> Avalon_FIR_0:avs_s0_write
	signal mm_interconnect_0_avalon_fir_0_s0_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_0:Avalon_FIR_0_s0_writedata -> Avalon_FIR_0:avs_s0_writedata
	signal mm_interconnect_0_onchip_memory_s1_chipselect            : std_logic;                     -- mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	signal mm_interconnect_0_onchip_memory_s1_readdata              : std_logic_vector(31 downto 0); -- onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	signal mm_interconnect_0_onchip_memory_s1_address               : std_logic_vector(9 downto 0);  -- mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	signal mm_interconnect_0_onchip_memory_s1_byteenable            : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	signal mm_interconnect_0_onchip_memory_s1_write                 : std_logic;                     -- mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	signal mm_interconnect_0_onchip_memory_s1_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	signal mm_interconnect_0_onchip_memory_s1_clken                 : std_logic;                     -- mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	signal mm_interconnect_0_jtag_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_avalon_jtag_slave_chipselect -> jtag:av_chipselect
	signal mm_interconnect_0_jtag_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag:av_readdata -> mm_interconnect_0:jtag_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag:av_waitrequest -> mm_interconnect_0:jtag_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_avalon_jtag_slave_address -> jtag:av_address
	signal mm_interconnect_0_jtag_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_avalon_jtag_slave_read -> mm_interconnect_0_jtag_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_avalon_jtag_slave_write -> mm_interconnect_0_jtag_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_avalon_jtag_slave_writedata -> jtag:av_writedata
	signal irq_mapper_receiver0_irq                                 : std_logic;                     -- jtag:av_irq -> irq_mapper:receiver0_irq
	signal nios_irq_irq                                             : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios:irq
	signal rst_controller_reset_out_reset                           : std_logic;                     -- rst_controller:reset_out -> [audio_config:reset, irq_mapper:reset, mm_interconnect_0:nios_reset_reset_bridge_in_reset_reset, onchip_memory:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                       : std_logic;                     -- rst_controller:reset_req -> [nios:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]
	signal reset_reset_n_ports_inv                                  : std_logic;                     -- reset_reset_n:inv -> [audio_pll:ref_reset_reset, rst_controller:reset_in0]
	signal mm_interconnect_0_jtag_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_avalon_jtag_slave_read:inv -> jtag:av_read_n
	signal mm_interconnect_0_jtag_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_avalon_jtag_slave_write:inv -> jtag:av_write_n
	signal rst_controller_reset_out_reset_ports_inv                 : std_logic;                     -- rst_controller_reset_out_reset:inv -> [AudioCodecAvalon_0:rsi_reset_n, Avalon_FIR_0:rsi_reset_n, jtag:rst_n, nios:reset_n]

begin

	audiocodecavalon_0 : component AudioCodecAvalon
		generic map (
			gDataWidth    => 24,
			gDataWidthLen => 5
		)
		port map (
			csi_clk         => clk_clk,                                      --        clock.clk
			rsi_reset_n     => rst_controller_reset_out_reset_ports_inv,     --        reset.reset_n
			AUD_ADCDAT      => i2s_adcdat,                                   --  conduit_end.adcdat
			AUD_ADCLRCK     => i2s_adclrck,                                  --             .adclrck
			AUD_BCLK        => i2s_bclk,                                     --             .bclk
			AUD_DACDAT      => i2s_dacdat,                                   --             .dacdat
			AUD_DACLRCK     => i2s_daclrck,                                  --             .daclrck
			asi_left_data   => avalon_fir_0_avalon_streaming_source_0_data,  --    left_sink.data
			asi_left_valid  => avalon_fir_0_avalon_streaming_source_0_valid, --             .valid
			asi_right_data  => audiocodecavalon_0_right_source_data,         --   right_sink.data
			asi_right_valid => audiocodecavalon_0_right_source_valid,        --             .valid
			aso_left_data   => audiocodecavalon_0_left_source_data,          --  left_source.data
			aso_left_valid  => audiocodecavalon_0_left_source_valid,         --             .valid
			aso_right_data  => audiocodecavalon_0_right_source_data,         -- right_source.data
			aso_right_valid => audiocodecavalon_0_right_source_valid         --             .valid
		);

	avalon_fir_0 : component FIR
		generic map (
			gDataWidth      => 24,
			gNrAddressLines => 4
		)
		port map (
			csi_clk          => clk_clk,                                      --                     clock.clk
			rsi_reset_n      => rst_controller_reset_out_reset_ports_inv,     --                     reset.reset_n
			avs_s0_address   => mm_interconnect_0_avalon_fir_0_s0_address,    --                        s0.address
			avs_s0_write     => mm_interconnect_0_avalon_fir_0_s0_write,      --                          .write
			avs_s0_writedata => mm_interconnect_0_avalon_fir_0_s0_writedata,  --                          .writedata
			avs_s0_read      => mm_interconnect_0_avalon_fir_0_s0_read,       --                          .read
			avs_s0_readdata  => mm_interconnect_0_avalon_fir_0_s0_readdata,   --                          .readdata
			asi_valid        => audiocodecavalon_0_left_source_valid,         --   avalon_streaming_sink_0.valid
			asi_data         => audiocodecavalon_0_left_source_data,          --                          .data
			aso_valid        => avalon_fir_0_avalon_streaming_source_0_valid, -- avalon_streaming_source_0.valid
			aso_data         => avalon_fir_0_avalon_streaming_source_0_data   --                          .data
		);

	audio_config : component Audio_audio_config
		port map (
			clk         => clk_clk,                        --                    clk.clk
			reset       => rst_controller_reset_out_reset, --                  reset.reset
			address     => open,                           -- avalon_av_config_slave.address
			byteenable  => open,                           --                       .byteenable
			read        => open,                           --                       .read
			write       => open,                           --                       .write
			writedata   => open,                           --                       .writedata
			readdata    => open,                           --                       .readdata
			waitrequest => open,                           --                       .waitrequest
			I2C_SDAT    => i2c_SDAT,                       --     external_interface.export
			I2C_SCLK    => i2c_SCLK                        --                       .export
		);

	audio_pll : component Audio_audio_pll
		port map (
			ref_clk_clk        => clk_clk,                 --      ref_clk.clk
			ref_reset_reset    => reset_reset_n_ports_inv, --    ref_reset.reset
			audio_clk_clk      => audio_clk_clk,           --    audio_clk.clk
			reset_source_reset => open                     -- reset_source.reset
		);

	jtag : component Audio_jtag
		port map (
			clk            => clk_clk,                                                  --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                 --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                  --               irq.irq
		);

	nios : component Audio_nios
		port map (
			clk                                 => clk_clk,                                            --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,           --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                 --                          .reset_req
			d_address                           => nios_data_master_address,                           --               data_master.address
			d_byteenable                        => nios_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios_data_master_read,                              --                          .read
			d_readdata                          => nios_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios_data_master_write,                             --                          .write
			d_writedata                         => nios_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios_instruction_master_read,                       --                          .read
			i_readdata                          => nios_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => open,                                               --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                -- custom_instruction_master.readra
		);

	onchip_memory : component Audio_onchip_memory
		port map (
			clk        => clk_clk,                                       --   clk1.clk
			address    => mm_interconnect_0_onchip_memory_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,            --       .reset_req
			freeze     => '0'                                            -- (terminated)
		);

	mm_interconnect_0 : component Audio_mm_interconnect_0
		port map (
			clk_clk_clk                            => clk_clk,                                              --                          clk_clk.clk
			nios_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                       -- nios_reset_reset_bridge_in_reset.reset
			nios_data_master_address               => nios_data_master_address,                             --                 nios_data_master.address
			nios_data_master_waitrequest           => nios_data_master_waitrequest,                         --                                 .waitrequest
			nios_data_master_byteenable            => nios_data_master_byteenable,                          --                                 .byteenable
			nios_data_master_read                  => nios_data_master_read,                                --                                 .read
			nios_data_master_readdata              => nios_data_master_readdata,                            --                                 .readdata
			nios_data_master_write                 => nios_data_master_write,                               --                                 .write
			nios_data_master_writedata             => nios_data_master_writedata,                           --                                 .writedata
			nios_data_master_debugaccess           => nios_data_master_debugaccess,                         --                                 .debugaccess
			nios_instruction_master_address        => nios_instruction_master_address,                      --          nios_instruction_master.address
			nios_instruction_master_waitrequest    => nios_instruction_master_waitrequest,                  --                                 .waitrequest
			nios_instruction_master_read           => nios_instruction_master_read,                         --                                 .read
			nios_instruction_master_readdata       => nios_instruction_master_readdata,                     --                                 .readdata
			Avalon_FIR_0_s0_address                => mm_interconnect_0_avalon_fir_0_s0_address,            --                  Avalon_FIR_0_s0.address
			Avalon_FIR_0_s0_write                  => mm_interconnect_0_avalon_fir_0_s0_write,              --                                 .write
			Avalon_FIR_0_s0_read                   => mm_interconnect_0_avalon_fir_0_s0_read,               --                                 .read
			Avalon_FIR_0_s0_readdata               => mm_interconnect_0_avalon_fir_0_s0_readdata,           --                                 .readdata
			Avalon_FIR_0_s0_writedata              => mm_interconnect_0_avalon_fir_0_s0_writedata,          --                                 .writedata
			jtag_avalon_jtag_slave_address         => mm_interconnect_0_jtag_avalon_jtag_slave_address,     --           jtag_avalon_jtag_slave.address
			jtag_avalon_jtag_slave_write           => mm_interconnect_0_jtag_avalon_jtag_slave_write,       --                                 .write
			jtag_avalon_jtag_slave_read            => mm_interconnect_0_jtag_avalon_jtag_slave_read,        --                                 .read
			jtag_avalon_jtag_slave_readdata        => mm_interconnect_0_jtag_avalon_jtag_slave_readdata,    --                                 .readdata
			jtag_avalon_jtag_slave_writedata       => mm_interconnect_0_jtag_avalon_jtag_slave_writedata,   --                                 .writedata
			jtag_avalon_jtag_slave_waitrequest     => mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest, --                                 .waitrequest
			jtag_avalon_jtag_slave_chipselect      => mm_interconnect_0_jtag_avalon_jtag_slave_chipselect,  --                                 .chipselect
			nios_debug_mem_slave_address           => mm_interconnect_0_nios_debug_mem_slave_address,       --             nios_debug_mem_slave.address
			nios_debug_mem_slave_write             => mm_interconnect_0_nios_debug_mem_slave_write,         --                                 .write
			nios_debug_mem_slave_read              => mm_interconnect_0_nios_debug_mem_slave_read,          --                                 .read
			nios_debug_mem_slave_readdata          => mm_interconnect_0_nios_debug_mem_slave_readdata,      --                                 .readdata
			nios_debug_mem_slave_writedata         => mm_interconnect_0_nios_debug_mem_slave_writedata,     --                                 .writedata
			nios_debug_mem_slave_byteenable        => mm_interconnect_0_nios_debug_mem_slave_byteenable,    --                                 .byteenable
			nios_debug_mem_slave_waitrequest       => mm_interconnect_0_nios_debug_mem_slave_waitrequest,   --                                 .waitrequest
			nios_debug_mem_slave_debugaccess       => mm_interconnect_0_nios_debug_mem_slave_debugaccess,   --                                 .debugaccess
			onchip_memory_s1_address               => mm_interconnect_0_onchip_memory_s1_address,           --                 onchip_memory_s1.address
			onchip_memory_s1_write                 => mm_interconnect_0_onchip_memory_s1_write,             --                                 .write
			onchip_memory_s1_readdata              => mm_interconnect_0_onchip_memory_s1_readdata,          --                                 .readdata
			onchip_memory_s1_writedata             => mm_interconnect_0_onchip_memory_s1_writedata,         --                                 .writedata
			onchip_memory_s1_byteenable            => mm_interconnect_0_onchip_memory_s1_byteenable,        --                                 .byteenable
			onchip_memory_s1_chipselect            => mm_interconnect_0_onchip_memory_s1_chipselect,        --                                 .chipselect
			onchip_memory_s1_clken                 => mm_interconnect_0_onchip_memory_s1_clken              --                                 .clken
		);

	irq_mapper : component Audio_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			sender_irq    => nios_irq_irq                    --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_avalon_jtag_slave_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of Audio
