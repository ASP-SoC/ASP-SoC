-- AudioSubSystem.vhd

-- Generated using ACDS version 16.1 196

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity AudioSubSystem is
	port (
		clk_clk       : in std_logic := '0'; --   clk.clk
		reset_reset_n : in std_logic := '0'  -- reset.reset_n
	);
end entity AudioSubSystem;

architecture rtl of AudioSubSystem is
	component AudioAvalonStream is
		port (
			clk                            : in  std_logic                     := 'X';             -- clk
			reset                          : in  std_logic                     := 'X';             -- reset_n
			from_audio_left_channel_data   : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			from_audio_left_channel_ready  : out std_logic;                                        -- ready
			from_audio_left_channel_valid  : in  std_logic                     := 'X';             -- valid
			from_audio_right_channel_data  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			from_audio_right_channel_ready : out std_logic;                                        -- ready
			from_audio_right_channel_valid : in  std_logic                     := 'X';             -- valid
			to_audio_left_channel_data     : out std_logic_vector(23 downto 0);                    -- data
			to_audio_left_channel_ready    : in  std_logic                     := 'X';             -- ready
			to_audio_left_channel_valid    : out std_logic;                                        -- valid
			to_audio_right_channel_data    : out std_logic_vector(23 downto 0);                    -- data
			to_audio_right_channel_ready   : in  std_logic                     := 'X';             -- ready
			to_audio_right_channel_valid   : out std_logic;                                        -- valid
			audio_sink_data                : in  std_logic_vector(47 downto 0) := (others => 'X'); -- data
			audio_sink_ready               : out std_logic;                                        -- ready
			audio_sink_valid               : in  std_logic                     := 'X';             -- valid
			audio_source_data              : out std_logic_vector(47 downto 0);                    -- data
			audio_source_valid             : out std_logic;                                        -- valid
			audio_source_ready             : in  std_logic                     := 'X'              -- ready
		);
	end component AudioAvalonStream;

	component AudioSubSystem_audio is
		port (
			clk                          : in  std_logic                     := 'X';             -- clk
			reset                        : in  std_logic                     := 'X';             -- reset
			from_adc_left_channel_ready  : in  std_logic                     := 'X';             -- ready
			from_adc_left_channel_data   : out std_logic_vector(23 downto 0);                    -- data
			from_adc_left_channel_valid  : out std_logic;                                        -- valid
			from_adc_right_channel_ready : in  std_logic                     := 'X';             -- ready
			from_adc_right_channel_data  : out std_logic_vector(23 downto 0);                    -- data
			from_adc_right_channel_valid : out std_logic;                                        -- valid
			to_dac_left_channel_data     : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			to_dac_left_channel_valid    : in  std_logic                     := 'X';             -- valid
			to_dac_left_channel_ready    : out std_logic;                                        -- ready
			to_dac_right_channel_data    : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			to_dac_right_channel_valid   : in  std_logic                     := 'X';             -- valid
			to_dac_right_channel_ready   : out std_logic;                                        -- ready
			AUD_ADCDAT                   : in  std_logic                     := 'X';             -- export
			AUD_ADCLRCK                  : in  std_logic                     := 'X';             -- export
			AUD_BCLK                     : in  std_logic                     := 'X';             -- export
			AUD_DACDAT                   : out std_logic;                                        -- export
			AUD_DACLRCK                  : in  std_logic                     := 'X'              -- export
		);
	end component AudioSubSystem_audio;

	component AudioSubSystem_audio_config is
		port (
			clk         : in    std_logic                     := 'X';             -- clk
			reset       : in    std_logic                     := 'X';             -- reset
			address     : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable  : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			read        : in    std_logic                     := 'X';             -- read
			write       : in    std_logic                     := 'X';             -- write
			writedata   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata    : out   std_logic_vector(31 downto 0);                    -- readdata
			waitrequest : out   std_logic;                                        -- waitrequest
			I2C_SDAT    : inout std_logic                     := 'X';             -- export
			I2C_SCLK    : out   std_logic                                         -- export
		);
	end component AudioSubSystem_audio_config;

	component AudioSubSystem_audio_pll is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			audio_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component AudioSubSystem_audio_pll;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal audioavalonstream_0_audio_left_channel_source_valid  : std_logic;                     -- AudioAvalonStream_0:to_audio_left_channel_valid -> audio:to_dac_left_channel_valid
	signal audioavalonstream_0_audio_left_channel_source_data   : std_logic_vector(23 downto 0); -- AudioAvalonStream_0:to_audio_left_channel_data -> audio:to_dac_left_channel_data
	signal audioavalonstream_0_audio_left_channel_source_ready  : std_logic;                     -- audio:to_dac_left_channel_ready -> AudioAvalonStream_0:to_audio_left_channel_ready
	signal audioavalonstream_0_audio_right_channel_source_valid : std_logic;                     -- AudioAvalonStream_0:to_audio_right_channel_valid -> audio:to_dac_right_channel_valid
	signal audioavalonstream_0_audio_right_channel_source_data  : std_logic_vector(23 downto 0); -- AudioAvalonStream_0:to_audio_right_channel_data -> audio:to_dac_right_channel_data
	signal audioavalonstream_0_audio_right_channel_source_ready : std_logic;                     -- audio:to_dac_right_channel_ready -> AudioAvalonStream_0:to_audio_right_channel_ready
	signal audioavalonstream_0_avalon_audio_source_valid        : std_logic;                     -- AudioAvalonStream_0:audio_source_valid -> AudioAvalonStream_0:audio_sink_valid
	signal audioavalonstream_0_avalon_audio_source_data         : std_logic_vector(47 downto 0); -- AudioAvalonStream_0:audio_source_data -> AudioAvalonStream_0:audio_sink_data
	signal audioavalonstream_0_avalon_audio_source_ready        : std_logic;                     -- AudioAvalonStream_0:audio_sink_ready -> AudioAvalonStream_0:audio_source_ready
	signal audio_avalon_left_channel_source_valid               : std_logic;                     -- audio:from_adc_left_channel_valid -> AudioAvalonStream_0:from_audio_left_channel_valid
	signal audio_avalon_left_channel_source_data                : std_logic_vector(23 downto 0); -- audio:from_adc_left_channel_data -> AudioAvalonStream_0:from_audio_left_channel_data
	signal audio_avalon_left_channel_source_ready               : std_logic;                     -- AudioAvalonStream_0:from_audio_left_channel_ready -> audio:from_adc_left_channel_ready
	signal audio_avalon_right_channel_source_valid              : std_logic;                     -- audio:from_adc_right_channel_valid -> AudioAvalonStream_0:from_audio_right_channel_valid
	signal audio_avalon_right_channel_source_data               : std_logic_vector(23 downto 0); -- audio:from_adc_right_channel_data -> AudioAvalonStream_0:from_audio_right_channel_data
	signal audio_avalon_right_channel_source_ready              : std_logic;                     -- AudioAvalonStream_0:from_audio_right_channel_ready -> audio:from_adc_right_channel_ready
	signal audio_pll_audio_clk_clk                              : std_logic;                     -- audio_pll:audio_clk_clk -> [AudioAvalonStream_0:clk, audio:clk, rst_controller:clk]
	signal rst_controller_reset_out_reset                       : std_logic;                     -- rst_controller:reset_out -> [audio:reset, rst_controller_reset_out_reset:in]
	signal audio_pll_reset_source_reset                         : std_logic;                     -- audio_pll:reset_source_reset -> rst_controller:reset_in0
	signal rst_controller_001_reset_out_reset                   : std_logic;                     -- rst_controller_001:reset_out -> audio_config:reset
	signal reset_reset_n_ports_inv                              : std_logic;                     -- reset_reset_n:inv -> [audio_pll:ref_reset_reset, rst_controller_001:reset_in0]
	signal rst_controller_reset_out_reset_ports_inv             : std_logic;                     -- rst_controller_reset_out_reset:inv -> AudioAvalonStream_0:reset

begin

	audioavalonstream_0 : component AudioAvalonStream
		port map (
			clk                            => audio_pll_audio_clk_clk,                              --                      clock.clk
			reset                          => rst_controller_reset_out_reset_ports_inv,             --                      reset.reset_n
			from_audio_left_channel_data   => audio_avalon_left_channel_source_data,                --    audio_left_channel_sink.data
			from_audio_left_channel_ready  => audio_avalon_left_channel_source_ready,               --                           .ready
			from_audio_left_channel_valid  => audio_avalon_left_channel_source_valid,               --                           .valid
			from_audio_right_channel_data  => audio_avalon_right_channel_source_data,               --   audio_right_channel_sink.data
			from_audio_right_channel_ready => audio_avalon_right_channel_source_ready,              --                           .ready
			from_audio_right_channel_valid => audio_avalon_right_channel_source_valid,              --                           .valid
			to_audio_left_channel_data     => audioavalonstream_0_audio_left_channel_source_data,   --  audio_left_channel_source.data
			to_audio_left_channel_ready    => audioavalonstream_0_audio_left_channel_source_ready,  --                           .ready
			to_audio_left_channel_valid    => audioavalonstream_0_audio_left_channel_source_valid,  --                           .valid
			to_audio_right_channel_data    => audioavalonstream_0_audio_right_channel_source_data,  -- audio_right_channel_source.data
			to_audio_right_channel_ready   => audioavalonstream_0_audio_right_channel_source_ready, --                           .ready
			to_audio_right_channel_valid   => audioavalonstream_0_audio_right_channel_source_valid, --                           .valid
			audio_sink_data                => audioavalonstream_0_avalon_audio_source_data,         --          avalon_audio_sink.data
			audio_sink_ready               => audioavalonstream_0_avalon_audio_source_ready,        --                           .ready
			audio_sink_valid               => audioavalonstream_0_avalon_audio_source_valid,        --                           .valid
			audio_source_data              => audioavalonstream_0_avalon_audio_source_data,         --        avalon_audio_source.data
			audio_source_valid             => audioavalonstream_0_avalon_audio_source_valid,        --                           .valid
			audio_source_ready             => audioavalonstream_0_avalon_audio_source_ready         --                           .ready
		);

	audio : component AudioSubSystem_audio
		port map (
			clk                          => audio_pll_audio_clk_clk,                              --                         clk.clk
			reset                        => rst_controller_reset_out_reset,                       --                       reset.reset
			from_adc_left_channel_ready  => audio_avalon_left_channel_source_ready,               --  avalon_left_channel_source.ready
			from_adc_left_channel_data   => audio_avalon_left_channel_source_data,                --                            .data
			from_adc_left_channel_valid  => audio_avalon_left_channel_source_valid,               --                            .valid
			from_adc_right_channel_ready => audio_avalon_right_channel_source_ready,              -- avalon_right_channel_source.ready
			from_adc_right_channel_data  => audio_avalon_right_channel_source_data,               --                            .data
			from_adc_right_channel_valid => audio_avalon_right_channel_source_valid,              --                            .valid
			to_dac_left_channel_data     => audioavalonstream_0_audio_left_channel_source_data,   --    avalon_left_channel_sink.data
			to_dac_left_channel_valid    => audioavalonstream_0_audio_left_channel_source_valid,  --                            .valid
			to_dac_left_channel_ready    => audioavalonstream_0_audio_left_channel_source_ready,  --                            .ready
			to_dac_right_channel_data    => audioavalonstream_0_audio_right_channel_source_data,  --   avalon_right_channel_sink.data
			to_dac_right_channel_valid   => audioavalonstream_0_audio_right_channel_source_valid, --                            .valid
			to_dac_right_channel_ready   => audioavalonstream_0_audio_right_channel_source_ready, --                            .ready
			AUD_ADCDAT                   => open,                                                 --          external_interface.export
			AUD_ADCLRCK                  => open,                                                 --                            .export
			AUD_BCLK                     => open,                                                 --                            .export
			AUD_DACDAT                   => open,                                                 --                            .export
			AUD_DACLRCK                  => open                                                  --                            .export
		);

	audio_config : component AudioSubSystem_audio_config
		port map (
			clk         => clk_clk,                            --                    clk.clk
			reset       => rst_controller_001_reset_out_reset, --                  reset.reset
			address     => open,                               -- avalon_av_config_slave.address
			byteenable  => open,                               --                       .byteenable
			read        => open,                               --                       .read
			write       => open,                               --                       .write
			writedata   => open,                               --                       .writedata
			readdata    => open,                               --                       .readdata
			waitrequest => open,                               --                       .waitrequest
			I2C_SDAT    => open,                               --     external_interface.export
			I2C_SCLK    => open                                --                       .export
		);

	audio_pll : component AudioSubSystem_audio_pll
		port map (
			ref_clk_clk        => clk_clk,                      --      ref_clk.clk
			ref_reset_reset    => reset_reset_n_ports_inv,      --    ref_reset.reset
			audio_clk_clk      => audio_pll_audio_clk_clk,      --    audio_clk.clk
			reset_source_reset => audio_pll_reset_source_reset  -- reset_source.reset
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => audio_pll_reset_source_reset,   -- reset_in0.reset
			clk            => audio_pll_audio_clk_clk,        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of AudioSubSystem
